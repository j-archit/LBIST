// ORA #2 - Comparator Module

module comp
#(parameter RC_BITS = 2)
(
    input [0 : RC_BITS - 1] rc_op,
    input [0 : RC_BITS - 1] ff_sig,
    output res
);
    
endmodule