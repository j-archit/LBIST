// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26
// Nfaults 902

module c880f (INC,END,clk,rst,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N72_t,N73_t,N74_t,N85_t,N86_t,N87_t,N88_t,N89_t,N90_t,N152_t,
     N259_t,N260_t,N267_t,N268_t;
wire N1_t0,N1_t1,N1_t2,N1_t3,N1_t4,N1_t5,N8_t0,N8_t1,N8_t2,
     N8_t3,N13_t0,N13_t1,N13_t2,N17_t0,N17_t1,N17_t2,N17_t3,N17_t4,N17_t5,
     N17_t6,N17_t7,N26_t0,N26_t1,N29_t0,N29_t1,N29_t2,N29_t3,N29_t4,N29_t5,
     N36_t0,N36_t1,N36_t2,N36_t3,N36_t4,N42_t0,N42_t1,N42_t2,N42_t3,N42_t4,
     N42_t5,N42_t6,N42_t7,N51_t0,N51_t1,N51_t2,N55_t0,N55_t1,N55_t2,N59_t0,
     N59_t1,N59_t2,N59_t3,N59_t4,N59_t5,N59_t6,N59_t7,N68_t0,N68_t1,N68_t2,
     N75_t0,N75_t1,N75_t2,N75_t3,N80_t0,N80_t1,N80_t2,N80_t3,N91_t0,N91_t1,
     N91_t2,N91_t3,N96_t0,N96_t1,N96_t2,N96_t3,N101_t0,N101_t1,N101_t2,N101_t3,
     N106_t0,N106_t1,N106_t2,N106_t3,N111_t0,N111_t1,N111_t2,N111_t3,N116_t0,N116_t1,
     N116_t2,N116_t3,N121_t0,N121_t1,N121_t2,N121_t3,N126_t0,N126_t1,N126_t2,N138_t0,
     N138_t1,N138_t2,N138_t3,N156_t0,N156_t1,N159_t0,N159_t1,N159_t2,N159_t3,N159_t4,
     N165_t0,N165_t1,N165_t2,N165_t3,N165_t4,N171_t0,N171_t1,N171_t2,N171_t3,N171_t4,
     N177_t0,N177_t1,N177_t2,N177_t3,N177_t4,N183_t0,N183_t1,N183_t2,N183_t3,N183_t4,
     N189_t0,N189_t1,N189_t2,N189_t3,N189_t4,N195_t0,N195_t1,N195_t2,N195_t3,N195_t4,
     N201_t0,N201_t1,N201_t2,N201_t3,N201_t4,N210_t0,N210_t1,N210_t2,N210_t3,N210_t4,
     N210_t5,N210_t6,N210_t7,N255_t0,N255_t1,N255_t2,N273_t0,N273_t1,N270_t0,N270_t1,
     N276_t0,N276_t1,N280_t0,N280_t1,N280_t2,N298_t0,N298_t1,N310_t0,N310_t1,N310_t2,
     N310_t3,N310_t4,N357_t0,N357_t1,N360_t0,N360_t1,N363_t0,N363_t1,N366_t0,N366_t1,
     N376_t0,N376_t1,N379_t0,N379_t1,N382_t0,N382_t1,N385_t0,N385_t1,N369_t0,N369_t1,
     N369_t2,N369_t3,N369_t4,N319_t0,N319_t1,N393_t0,N393_t1,N393_t2,N393_t3,N393_t4,
     N287_t0,N287_t1,N143_t0,N143_t1,N427_t0,N427_t1,N427_t2,N427_t3,N432_t0,N432_t1,
     N432_t2,N432_t3,N146_t0,N146_t1,N149_t0,N149_t1,N153_t0,N153_t1,N437_t0,N437_t1,
     N437_t2,N437_t3,N130_t0,N130_t1,N130_t2,N130_t3,N460_t0,N460_t1,N463_t0,N463_t1,
     N135_t0,N135_t1,N466_t0,N466_t1,N466_t2,N466_t3,N466_t4,N466_t5,N466_t6,N466_t7,
     N483_t0,N483_t1,N483_t2,N483_t3,N492_t0,N492_t1,N495_t0,N495_t1,N207_t0,N207_t1,
     N451_t0,N451_t1,N451_t2,N451_t3,N451_t4,N451_t5,N451_t6,N451_t7,N530_t0,N530_t1,
     N533_t0,N533_t1,N544_t0,N544_t1,N547_t0,N547_t1,N553_t0,N553_t1,N553_t2,N246_t0,
     N246_t1,N246_t2,N246_t3,N246_t4,N246_t5,N246_t6,N246_t7,N557_t0,N557_t1,N557_t2,
     N561_t0,N561_t1,N561_t2,N565_t0,N565_t1,N565_t2,N569_t0,N569_t1,N569_t2,N573_t0,
     N573_t1,N573_t2,N577_t0,N577_t1,N577_t2,N581_t0,N581_t1,N581_t2,N590_t0,N590_t1,
     N593_t0,N593_t1,N597_t0,N597_t1,N600_t0,N600_t1,N600_t2,N600_t3,N606_t0,N606_t1,
     N609_t0,N609_t1,N609_t2,N609_t3,N609_t4,N616_t0,N616_t1,N619_t0,N619_t1,N619_t2,
     N619_t3,N625_t0,N625_t1,N628_t0,N628_t1,N632_t0,N632_t1,N635_t0,N635_t1,N635_t2,
     N635_t3,N641_t0,N641_t1,N644_t0,N644_t1,N644_t2,N644_t3,N644_t4,N651_t0,N651_t1,
     N654_t0,N654_t1,N654_t2,N654_t3,N261_t0,N261_t1,N261_t2,N261_t3,N261_t4,N662_t0,
     N662_t1,N228_t0,N228_t1,N228_t2,N228_t3,N228_t4,N228_t5,N228_t6,N228_t7,N665_t0,
     N665_t1,N665_t2,N237_t0,N237_t1,N237_t2,N237_t3,N237_t4,N237_t5,N237_t6,N237_t7,
     N670_t0,N670_t1,N673_t0,N673_t1,N673_t2,N678_t0,N678_t1,N678_t2,N682_t0,N682_t1,
     N682_t2,N687_t0,N687_t1,N687_t2,N687_t3,N692_t0,N692_t1,N692_t2,N697_t0,N697_t1,
     N700_t0,N700_t1,N700_t2,N705_t0,N705_t1,N708_t0,N708_t1,N708_t2,N713_t0,N713_t1,
     N713_t2,N717_t0,N717_t1,N717_t2,N722_t0,N722_t1,N722_t2,N722_t3,N727_t0,N727_t1,
     N727_t2,N773_t0,N773_t1,N773_t2,N778_t0,N778_t1,N782_t0,N782_t1,N219_t0,N219_t1,
     N219_t2,N219_t3,N219_t4,N219_t5,N219_t6,N219_t7,N796_t0,N796_t1,N796_t2,N796_t3,
     N796_t4,N815_t0,N815_t1,N815_t2,N819_t0,N819_t1,N822_t0,N822_t1;
reg [450:0] FEN;
fim PI_N72( .fault(fault), .net(N72), .FEN(FEN[0]), .op(N72_t) );
fim PI_N73( .fault(fault), .net(N73), .FEN(FEN[1]), .op(N73_t) );
fim PI_N74( .fault(fault), .net(N74), .FEN(FEN[2]), .op(N74_t) );
fim PI_N85( .fault(fault), .net(N85), .FEN(FEN[3]), .op(N85_t) );
fim PI_N86( .fault(fault), .net(N86), .FEN(FEN[4]), .op(N86_t) );
fim PI_N87( .fault(fault), .net(N87), .FEN(FEN[5]), .op(N87_t) );
fim PI_N88( .fault(fault), .net(N88), .FEN(FEN[6]), .op(N88_t) );
fim PI_N89( .fault(fault), .net(N89), .FEN(FEN[7]), .op(N89_t) );
fim PI_N90( .fault(fault), .net(N90), .FEN(FEN[8]), .op(N90_t) );
fim PI_N152( .fault(fault), .net(N152), .FEN(FEN[9]), .op(N152_t) );
fim PI_N259( .fault(fault), .net(N259), .FEN(FEN[10]), .op(N259_t) );
fim PI_N260( .fault(fault), .net(N260), .FEN(FEN[11]), .op(N260_t) );
fim PI_N267( .fault(fault), .net(N267), .FEN(FEN[12]), .op(N267_t) );
fim PI_N268( .fault(fault), .net(N268), .FEN(FEN[13]), .op(N268_t) );
fim FAN_N1_0 ( .fault(fault), .net(N1), .FEN(FEN[14]), .op(N1_t0) );
fim FAN_N1_1 ( .fault(fault), .net(N1), .FEN(FEN[15]), .op(N1_t1) );
fim FAN_N1_2 ( .fault(fault), .net(N1), .FEN(FEN[16]), .op(N1_t2) );
fim FAN_N1_3 ( .fault(fault), .net(N1), .FEN(FEN[17]), .op(N1_t3) );
fim FAN_N1_4 ( .fault(fault), .net(N1), .FEN(FEN[18]), .op(N1_t4) );
fim FAN_N1_5 ( .fault(fault), .net(N1), .FEN(FEN[19]), .op(N1_t5) );
fim FAN_N8_0 ( .fault(fault), .net(N8), .FEN(FEN[20]), .op(N8_t0) );
fim FAN_N8_1 ( .fault(fault), .net(N8), .FEN(FEN[21]), .op(N8_t1) );
fim FAN_N8_2 ( .fault(fault), .net(N8), .FEN(FEN[22]), .op(N8_t2) );
fim FAN_N8_3 ( .fault(fault), .net(N8), .FEN(FEN[23]), .op(N8_t3) );
fim FAN_N13_0 ( .fault(fault), .net(N13), .FEN(FEN[24]), .op(N13_t0) );
fim FAN_N13_1 ( .fault(fault), .net(N13), .FEN(FEN[25]), .op(N13_t1) );
fim FAN_N13_2 ( .fault(fault), .net(N13), .FEN(FEN[26]), .op(N13_t2) );
fim FAN_N17_0 ( .fault(fault), .net(N17), .FEN(FEN[27]), .op(N17_t0) );
fim FAN_N17_1 ( .fault(fault), .net(N17), .FEN(FEN[28]), .op(N17_t1) );
fim FAN_N17_2 ( .fault(fault), .net(N17), .FEN(FEN[29]), .op(N17_t2) );
fim FAN_N17_3 ( .fault(fault), .net(N17), .FEN(FEN[30]), .op(N17_t3) );
fim FAN_N17_4 ( .fault(fault), .net(N17), .FEN(FEN[31]), .op(N17_t4) );
fim FAN_N17_5 ( .fault(fault), .net(N17), .FEN(FEN[32]), .op(N17_t5) );
fim FAN_N17_6 ( .fault(fault), .net(N17), .FEN(FEN[33]), .op(N17_t6) );
fim FAN_N17_7 ( .fault(fault), .net(N17), .FEN(FEN[34]), .op(N17_t7) );
fim FAN_N26_0 ( .fault(fault), .net(N26), .FEN(FEN[35]), .op(N26_t0) );
fim FAN_N26_1 ( .fault(fault), .net(N26), .FEN(FEN[36]), .op(N26_t1) );
fim FAN_N29_0 ( .fault(fault), .net(N29), .FEN(FEN[37]), .op(N29_t0) );
fim FAN_N29_1 ( .fault(fault), .net(N29), .FEN(FEN[38]), .op(N29_t1) );
fim FAN_N29_2 ( .fault(fault), .net(N29), .FEN(FEN[39]), .op(N29_t2) );
fim FAN_N29_3 ( .fault(fault), .net(N29), .FEN(FEN[40]), .op(N29_t3) );
fim FAN_N29_4 ( .fault(fault), .net(N29), .FEN(FEN[41]), .op(N29_t4) );
fim FAN_N29_5 ( .fault(fault), .net(N29), .FEN(FEN[42]), .op(N29_t5) );
fim FAN_N36_0 ( .fault(fault), .net(N36), .FEN(FEN[43]), .op(N36_t0) );
fim FAN_N36_1 ( .fault(fault), .net(N36), .FEN(FEN[44]), .op(N36_t1) );
fim FAN_N36_2 ( .fault(fault), .net(N36), .FEN(FEN[45]), .op(N36_t2) );
fim FAN_N36_3 ( .fault(fault), .net(N36), .FEN(FEN[46]), .op(N36_t3) );
fim FAN_N36_4 ( .fault(fault), .net(N36), .FEN(FEN[47]), .op(N36_t4) );
fim FAN_N42_0 ( .fault(fault), .net(N42), .FEN(FEN[48]), .op(N42_t0) );
fim FAN_N42_1 ( .fault(fault), .net(N42), .FEN(FEN[49]), .op(N42_t1) );
fim FAN_N42_2 ( .fault(fault), .net(N42), .FEN(FEN[50]), .op(N42_t2) );
fim FAN_N42_3 ( .fault(fault), .net(N42), .FEN(FEN[51]), .op(N42_t3) );
fim FAN_N42_4 ( .fault(fault), .net(N42), .FEN(FEN[52]), .op(N42_t4) );
fim FAN_N42_5 ( .fault(fault), .net(N42), .FEN(FEN[53]), .op(N42_t5) );
fim FAN_N42_6 ( .fault(fault), .net(N42), .FEN(FEN[54]), .op(N42_t6) );
fim FAN_N42_7 ( .fault(fault), .net(N42), .FEN(FEN[55]), .op(N42_t7) );
fim FAN_N51_0 ( .fault(fault), .net(N51), .FEN(FEN[56]), .op(N51_t0) );
fim FAN_N51_1 ( .fault(fault), .net(N51), .FEN(FEN[57]), .op(N51_t1) );
fim FAN_N51_2 ( .fault(fault), .net(N51), .FEN(FEN[58]), .op(N51_t2) );
fim FAN_N55_0 ( .fault(fault), .net(N55), .FEN(FEN[59]), .op(N55_t0) );
fim FAN_N55_1 ( .fault(fault), .net(N55), .FEN(FEN[60]), .op(N55_t1) );
fim FAN_N55_2 ( .fault(fault), .net(N55), .FEN(FEN[61]), .op(N55_t2) );
fim FAN_N59_0 ( .fault(fault), .net(N59), .FEN(FEN[62]), .op(N59_t0) );
fim FAN_N59_1 ( .fault(fault), .net(N59), .FEN(FEN[63]), .op(N59_t1) );
fim FAN_N59_2 ( .fault(fault), .net(N59), .FEN(FEN[64]), .op(N59_t2) );
fim FAN_N59_3 ( .fault(fault), .net(N59), .FEN(FEN[65]), .op(N59_t3) );
fim FAN_N59_4 ( .fault(fault), .net(N59), .FEN(FEN[66]), .op(N59_t4) );
fim FAN_N59_5 ( .fault(fault), .net(N59), .FEN(FEN[67]), .op(N59_t5) );
fim FAN_N59_6 ( .fault(fault), .net(N59), .FEN(FEN[68]), .op(N59_t6) );
fim FAN_N59_7 ( .fault(fault), .net(N59), .FEN(FEN[69]), .op(N59_t7) );
fim FAN_N68_0 ( .fault(fault), .net(N68), .FEN(FEN[70]), .op(N68_t0) );
fim FAN_N68_1 ( .fault(fault), .net(N68), .FEN(FEN[71]), .op(N68_t1) );
fim FAN_N68_2 ( .fault(fault), .net(N68), .FEN(FEN[72]), .op(N68_t2) );
fim FAN_N75_0 ( .fault(fault), .net(N75), .FEN(FEN[73]), .op(N75_t0) );
fim FAN_N75_1 ( .fault(fault), .net(N75), .FEN(FEN[74]), .op(N75_t1) );
fim FAN_N75_2 ( .fault(fault), .net(N75), .FEN(FEN[75]), .op(N75_t2) );
fim FAN_N75_3 ( .fault(fault), .net(N75), .FEN(FEN[76]), .op(N75_t3) );
fim FAN_N80_0 ( .fault(fault), .net(N80), .FEN(FEN[77]), .op(N80_t0) );
fim FAN_N80_1 ( .fault(fault), .net(N80), .FEN(FEN[78]), .op(N80_t1) );
fim FAN_N80_2 ( .fault(fault), .net(N80), .FEN(FEN[79]), .op(N80_t2) );
fim FAN_N80_3 ( .fault(fault), .net(N80), .FEN(FEN[80]), .op(N80_t3) );
fim FAN_N91_0 ( .fault(fault), .net(N91), .FEN(FEN[81]), .op(N91_t0) );
fim FAN_N91_1 ( .fault(fault), .net(N91), .FEN(FEN[82]), .op(N91_t1) );
fim FAN_N91_2 ( .fault(fault), .net(N91), .FEN(FEN[83]), .op(N91_t2) );
fim FAN_N91_3 ( .fault(fault), .net(N91), .FEN(FEN[84]), .op(N91_t3) );
fim FAN_N96_0 ( .fault(fault), .net(N96), .FEN(FEN[85]), .op(N96_t0) );
fim FAN_N96_1 ( .fault(fault), .net(N96), .FEN(FEN[86]), .op(N96_t1) );
fim FAN_N96_2 ( .fault(fault), .net(N96), .FEN(FEN[87]), .op(N96_t2) );
fim FAN_N96_3 ( .fault(fault), .net(N96), .FEN(FEN[88]), .op(N96_t3) );
fim FAN_N101_0 ( .fault(fault), .net(N101), .FEN(FEN[89]), .op(N101_t0) );
fim FAN_N101_1 ( .fault(fault), .net(N101), .FEN(FEN[90]), .op(N101_t1) );
fim FAN_N101_2 ( .fault(fault), .net(N101), .FEN(FEN[91]), .op(N101_t2) );
fim FAN_N101_3 ( .fault(fault), .net(N101), .FEN(FEN[92]), .op(N101_t3) );
fim FAN_N106_0 ( .fault(fault), .net(N106), .FEN(FEN[93]), .op(N106_t0) );
fim FAN_N106_1 ( .fault(fault), .net(N106), .FEN(FEN[94]), .op(N106_t1) );
fim FAN_N106_2 ( .fault(fault), .net(N106), .FEN(FEN[95]), .op(N106_t2) );
fim FAN_N106_3 ( .fault(fault), .net(N106), .FEN(FEN[96]), .op(N106_t3) );
fim FAN_N111_0 ( .fault(fault), .net(N111), .FEN(FEN[97]), .op(N111_t0) );
fim FAN_N111_1 ( .fault(fault), .net(N111), .FEN(FEN[98]), .op(N111_t1) );
fim FAN_N111_2 ( .fault(fault), .net(N111), .FEN(FEN[99]), .op(N111_t2) );
fim FAN_N111_3 ( .fault(fault), .net(N111), .FEN(FEN[100]), .op(N111_t3) );
fim FAN_N116_0 ( .fault(fault), .net(N116), .FEN(FEN[101]), .op(N116_t0) );
fim FAN_N116_1 ( .fault(fault), .net(N116), .FEN(FEN[102]), .op(N116_t1) );
fim FAN_N116_2 ( .fault(fault), .net(N116), .FEN(FEN[103]), .op(N116_t2) );
fim FAN_N116_3 ( .fault(fault), .net(N116), .FEN(FEN[104]), .op(N116_t3) );
fim FAN_N121_0 ( .fault(fault), .net(N121), .FEN(FEN[105]), .op(N121_t0) );
fim FAN_N121_1 ( .fault(fault), .net(N121), .FEN(FEN[106]), .op(N121_t1) );
fim FAN_N121_2 ( .fault(fault), .net(N121), .FEN(FEN[107]), .op(N121_t2) );
fim FAN_N121_3 ( .fault(fault), .net(N121), .FEN(FEN[108]), .op(N121_t3) );
fim FAN_N126_0 ( .fault(fault), .net(N126), .FEN(FEN[109]), .op(N126_t0) );
fim FAN_N126_1 ( .fault(fault), .net(N126), .FEN(FEN[110]), .op(N126_t1) );
fim FAN_N126_2 ( .fault(fault), .net(N126), .FEN(FEN[111]), .op(N126_t2) );
fim FAN_N138_0 ( .fault(fault), .net(N138), .FEN(FEN[112]), .op(N138_t0) );
fim FAN_N138_1 ( .fault(fault), .net(N138), .FEN(FEN[113]), .op(N138_t1) );
fim FAN_N138_2 ( .fault(fault), .net(N138), .FEN(FEN[114]), .op(N138_t2) );
fim FAN_N138_3 ( .fault(fault), .net(N138), .FEN(FEN[115]), .op(N138_t3) );
fim FAN_N156_0 ( .fault(fault), .net(N156), .FEN(FEN[116]), .op(N156_t0) );
fim FAN_N156_1 ( .fault(fault), .net(N156), .FEN(FEN[117]), .op(N156_t1) );
fim FAN_N159_0 ( .fault(fault), .net(N159), .FEN(FEN[118]), .op(N159_t0) );
fim FAN_N159_1 ( .fault(fault), .net(N159), .FEN(FEN[119]), .op(N159_t1) );
fim FAN_N159_2 ( .fault(fault), .net(N159), .FEN(FEN[120]), .op(N159_t2) );
fim FAN_N159_3 ( .fault(fault), .net(N159), .FEN(FEN[121]), .op(N159_t3) );
fim FAN_N159_4 ( .fault(fault), .net(N159), .FEN(FEN[122]), .op(N159_t4) );
fim FAN_N165_0 ( .fault(fault), .net(N165), .FEN(FEN[123]), .op(N165_t0) );
fim FAN_N165_1 ( .fault(fault), .net(N165), .FEN(FEN[124]), .op(N165_t1) );
fim FAN_N165_2 ( .fault(fault), .net(N165), .FEN(FEN[125]), .op(N165_t2) );
fim FAN_N165_3 ( .fault(fault), .net(N165), .FEN(FEN[126]), .op(N165_t3) );
fim FAN_N165_4 ( .fault(fault), .net(N165), .FEN(FEN[127]), .op(N165_t4) );
fim FAN_N171_0 ( .fault(fault), .net(N171), .FEN(FEN[128]), .op(N171_t0) );
fim FAN_N171_1 ( .fault(fault), .net(N171), .FEN(FEN[129]), .op(N171_t1) );
fim FAN_N171_2 ( .fault(fault), .net(N171), .FEN(FEN[130]), .op(N171_t2) );
fim FAN_N171_3 ( .fault(fault), .net(N171), .FEN(FEN[131]), .op(N171_t3) );
fim FAN_N171_4 ( .fault(fault), .net(N171), .FEN(FEN[132]), .op(N171_t4) );
fim FAN_N177_0 ( .fault(fault), .net(N177), .FEN(FEN[133]), .op(N177_t0) );
fim FAN_N177_1 ( .fault(fault), .net(N177), .FEN(FEN[134]), .op(N177_t1) );
fim FAN_N177_2 ( .fault(fault), .net(N177), .FEN(FEN[135]), .op(N177_t2) );
fim FAN_N177_3 ( .fault(fault), .net(N177), .FEN(FEN[136]), .op(N177_t3) );
fim FAN_N177_4 ( .fault(fault), .net(N177), .FEN(FEN[137]), .op(N177_t4) );
fim FAN_N183_0 ( .fault(fault), .net(N183), .FEN(FEN[138]), .op(N183_t0) );
fim FAN_N183_1 ( .fault(fault), .net(N183), .FEN(FEN[139]), .op(N183_t1) );
fim FAN_N183_2 ( .fault(fault), .net(N183), .FEN(FEN[140]), .op(N183_t2) );
fim FAN_N183_3 ( .fault(fault), .net(N183), .FEN(FEN[141]), .op(N183_t3) );
fim FAN_N183_4 ( .fault(fault), .net(N183), .FEN(FEN[142]), .op(N183_t4) );
fim FAN_N189_0 ( .fault(fault), .net(N189), .FEN(FEN[143]), .op(N189_t0) );
fim FAN_N189_1 ( .fault(fault), .net(N189), .FEN(FEN[144]), .op(N189_t1) );
fim FAN_N189_2 ( .fault(fault), .net(N189), .FEN(FEN[145]), .op(N189_t2) );
fim FAN_N189_3 ( .fault(fault), .net(N189), .FEN(FEN[146]), .op(N189_t3) );
fim FAN_N189_4 ( .fault(fault), .net(N189), .FEN(FEN[147]), .op(N189_t4) );
fim FAN_N195_0 ( .fault(fault), .net(N195), .FEN(FEN[148]), .op(N195_t0) );
fim FAN_N195_1 ( .fault(fault), .net(N195), .FEN(FEN[149]), .op(N195_t1) );
fim FAN_N195_2 ( .fault(fault), .net(N195), .FEN(FEN[150]), .op(N195_t2) );
fim FAN_N195_3 ( .fault(fault), .net(N195), .FEN(FEN[151]), .op(N195_t3) );
fim FAN_N195_4 ( .fault(fault), .net(N195), .FEN(FEN[152]), .op(N195_t4) );
fim FAN_N201_0 ( .fault(fault), .net(N201), .FEN(FEN[153]), .op(N201_t0) );
fim FAN_N201_1 ( .fault(fault), .net(N201), .FEN(FEN[154]), .op(N201_t1) );
fim FAN_N201_2 ( .fault(fault), .net(N201), .FEN(FEN[155]), .op(N201_t2) );
fim FAN_N201_3 ( .fault(fault), .net(N201), .FEN(FEN[156]), .op(N201_t3) );
fim FAN_N201_4 ( .fault(fault), .net(N201), .FEN(FEN[157]), .op(N201_t4) );
fim FAN_N210_0 ( .fault(fault), .net(N210), .FEN(FEN[158]), .op(N210_t0) );
fim FAN_N210_1 ( .fault(fault), .net(N210), .FEN(FEN[159]), .op(N210_t1) );
fim FAN_N210_2 ( .fault(fault), .net(N210), .FEN(FEN[160]), .op(N210_t2) );
fim FAN_N210_3 ( .fault(fault), .net(N210), .FEN(FEN[161]), .op(N210_t3) );
fim FAN_N210_4 ( .fault(fault), .net(N210), .FEN(FEN[162]), .op(N210_t4) );
fim FAN_N210_5 ( .fault(fault), .net(N210), .FEN(FEN[163]), .op(N210_t5) );
fim FAN_N210_6 ( .fault(fault), .net(N210), .FEN(FEN[164]), .op(N210_t6) );
fim FAN_N210_7 ( .fault(fault), .net(N210), .FEN(FEN[165]), .op(N210_t7) );
fim FAN_N255_0 ( .fault(fault), .net(N255), .FEN(FEN[166]), .op(N255_t0) );
fim FAN_N255_1 ( .fault(fault), .net(N255), .FEN(FEN[167]), .op(N255_t1) );
fim FAN_N255_2 ( .fault(fault), .net(N255), .FEN(FEN[168]), .op(N255_t2) );
fim FAN_N273_0 ( .fault(fault), .net(N273), .FEN(FEN[169]), .op(N273_t0) );
fim FAN_N273_1 ( .fault(fault), .net(N273), .FEN(FEN[170]), .op(N273_t1) );
fim FAN_N270_0 ( .fault(fault), .net(N270), .FEN(FEN[171]), .op(N270_t0) );
fim FAN_N270_1 ( .fault(fault), .net(N270), .FEN(FEN[172]), .op(N270_t1) );
fim FAN_N276_0 ( .fault(fault), .net(N276), .FEN(FEN[173]), .op(N276_t0) );
fim FAN_N276_1 ( .fault(fault), .net(N276), .FEN(FEN[174]), .op(N276_t1) );
fim FAN_N280_0 ( .fault(fault), .net(N280), .FEN(FEN[175]), .op(N280_t0) );
fim FAN_N280_1 ( .fault(fault), .net(N280), .FEN(FEN[176]), .op(N280_t1) );
fim FAN_N280_2 ( .fault(fault), .net(N280), .FEN(FEN[177]), .op(N280_t2) );
fim FAN_N298_0 ( .fault(fault), .net(N298), .FEN(FEN[178]), .op(N298_t0) );
fim FAN_N298_1 ( .fault(fault), .net(N298), .FEN(FEN[179]), .op(N298_t1) );
fim FAN_N310_0 ( .fault(fault), .net(N310), .FEN(FEN[180]), .op(N310_t0) );
fim FAN_N310_1 ( .fault(fault), .net(N310), .FEN(FEN[181]), .op(N310_t1) );
fim FAN_N310_2 ( .fault(fault), .net(N310), .FEN(FEN[182]), .op(N310_t2) );
fim FAN_N310_3 ( .fault(fault), .net(N310), .FEN(FEN[183]), .op(N310_t3) );
fim FAN_N310_4 ( .fault(fault), .net(N310), .FEN(FEN[184]), .op(N310_t4) );
fim FAN_N357_0 ( .fault(fault), .net(N357), .FEN(FEN[185]), .op(N357_t0) );
fim FAN_N357_1 ( .fault(fault), .net(N357), .FEN(FEN[186]), .op(N357_t1) );
fim FAN_N360_0 ( .fault(fault), .net(N360), .FEN(FEN[187]), .op(N360_t0) );
fim FAN_N360_1 ( .fault(fault), .net(N360), .FEN(FEN[188]), .op(N360_t1) );
fim FAN_N363_0 ( .fault(fault), .net(N363), .FEN(FEN[189]), .op(N363_t0) );
fim FAN_N363_1 ( .fault(fault), .net(N363), .FEN(FEN[190]), .op(N363_t1) );
fim FAN_N366_0 ( .fault(fault), .net(N366), .FEN(FEN[191]), .op(N366_t0) );
fim FAN_N366_1 ( .fault(fault), .net(N366), .FEN(FEN[192]), .op(N366_t1) );
fim FAN_N376_0 ( .fault(fault), .net(N376), .FEN(FEN[193]), .op(N376_t0) );
fim FAN_N376_1 ( .fault(fault), .net(N376), .FEN(FEN[194]), .op(N376_t1) );
fim FAN_N379_0 ( .fault(fault), .net(N379), .FEN(FEN[195]), .op(N379_t0) );
fim FAN_N379_1 ( .fault(fault), .net(N379), .FEN(FEN[196]), .op(N379_t1) );
fim FAN_N382_0 ( .fault(fault), .net(N382), .FEN(FEN[197]), .op(N382_t0) );
fim FAN_N382_1 ( .fault(fault), .net(N382), .FEN(FEN[198]), .op(N382_t1) );
fim FAN_N385_0 ( .fault(fault), .net(N385), .FEN(FEN[199]), .op(N385_t0) );
fim FAN_N385_1 ( .fault(fault), .net(N385), .FEN(FEN[200]), .op(N385_t1) );
fim FAN_N369_0 ( .fault(fault), .net(N369), .FEN(FEN[201]), .op(N369_t0) );
fim FAN_N369_1 ( .fault(fault), .net(N369), .FEN(FEN[202]), .op(N369_t1) );
fim FAN_N369_2 ( .fault(fault), .net(N369), .FEN(FEN[203]), .op(N369_t2) );
fim FAN_N369_3 ( .fault(fault), .net(N369), .FEN(FEN[204]), .op(N369_t3) );
fim FAN_N369_4 ( .fault(fault), .net(N369), .FEN(FEN[205]), .op(N369_t4) );
fim FAN_N319_0 ( .fault(fault), .net(N319), .FEN(FEN[206]), .op(N319_t0) );
fim FAN_N319_1 ( .fault(fault), .net(N319), .FEN(FEN[207]), .op(N319_t1) );
fim FAN_N393_0 ( .fault(fault), .net(N393), .FEN(FEN[208]), .op(N393_t0) );
fim FAN_N393_1 ( .fault(fault), .net(N393), .FEN(FEN[209]), .op(N393_t1) );
fim FAN_N393_2 ( .fault(fault), .net(N393), .FEN(FEN[210]), .op(N393_t2) );
fim FAN_N393_3 ( .fault(fault), .net(N393), .FEN(FEN[211]), .op(N393_t3) );
fim FAN_N393_4 ( .fault(fault), .net(N393), .FEN(FEN[212]), .op(N393_t4) );
fim FAN_N287_0 ( .fault(fault), .net(N287), .FEN(FEN[213]), .op(N287_t0) );
fim FAN_N287_1 ( .fault(fault), .net(N287), .FEN(FEN[214]), .op(N287_t1) );
fim FAN_N143_0 ( .fault(fault), .net(N143), .FEN(FEN[215]), .op(N143_t0) );
fim FAN_N143_1 ( .fault(fault), .net(N143), .FEN(FEN[216]), .op(N143_t1) );
fim FAN_N427_0 ( .fault(fault), .net(N427), .FEN(FEN[217]), .op(N427_t0) );
fim FAN_N427_1 ( .fault(fault), .net(N427), .FEN(FEN[218]), .op(N427_t1) );
fim FAN_N427_2 ( .fault(fault), .net(N427), .FEN(FEN[219]), .op(N427_t2) );
fim FAN_N427_3 ( .fault(fault), .net(N427), .FEN(FEN[220]), .op(N427_t3) );
fim FAN_N432_0 ( .fault(fault), .net(N432), .FEN(FEN[221]), .op(N432_t0) );
fim FAN_N432_1 ( .fault(fault), .net(N432), .FEN(FEN[222]), .op(N432_t1) );
fim FAN_N432_2 ( .fault(fault), .net(N432), .FEN(FEN[223]), .op(N432_t2) );
fim FAN_N432_3 ( .fault(fault), .net(N432), .FEN(FEN[224]), .op(N432_t3) );
fim FAN_N146_0 ( .fault(fault), .net(N146), .FEN(FEN[225]), .op(N146_t0) );
fim FAN_N146_1 ( .fault(fault), .net(N146), .FEN(FEN[226]), .op(N146_t1) );
fim FAN_N149_0 ( .fault(fault), .net(N149), .FEN(FEN[227]), .op(N149_t0) );
fim FAN_N149_1 ( .fault(fault), .net(N149), .FEN(FEN[228]), .op(N149_t1) );
fim FAN_N153_0 ( .fault(fault), .net(N153), .FEN(FEN[229]), .op(N153_t0) );
fim FAN_N153_1 ( .fault(fault), .net(N153), .FEN(FEN[230]), .op(N153_t1) );
fim FAN_N437_0 ( .fault(fault), .net(N437), .FEN(FEN[231]), .op(N437_t0) );
fim FAN_N437_1 ( .fault(fault), .net(N437), .FEN(FEN[232]), .op(N437_t1) );
fim FAN_N437_2 ( .fault(fault), .net(N437), .FEN(FEN[233]), .op(N437_t2) );
fim FAN_N437_3 ( .fault(fault), .net(N437), .FEN(FEN[234]), .op(N437_t3) );
fim FAN_N130_0 ( .fault(fault), .net(N130), .FEN(FEN[235]), .op(N130_t0) );
fim FAN_N130_1 ( .fault(fault), .net(N130), .FEN(FEN[236]), .op(N130_t1) );
fim FAN_N130_2 ( .fault(fault), .net(N130), .FEN(FEN[237]), .op(N130_t2) );
fim FAN_N130_3 ( .fault(fault), .net(N130), .FEN(FEN[238]), .op(N130_t3) );
fim FAN_N460_0 ( .fault(fault), .net(N460), .FEN(FEN[239]), .op(N460_t0) );
fim FAN_N460_1 ( .fault(fault), .net(N460), .FEN(FEN[240]), .op(N460_t1) );
fim FAN_N463_0 ( .fault(fault), .net(N463), .FEN(FEN[241]), .op(N463_t0) );
fim FAN_N463_1 ( .fault(fault), .net(N463), .FEN(FEN[242]), .op(N463_t1) );
fim FAN_N135_0 ( .fault(fault), .net(N135), .FEN(FEN[243]), .op(N135_t0) );
fim FAN_N135_1 ( .fault(fault), .net(N135), .FEN(FEN[244]), .op(N135_t1) );
fim FAN_N466_0 ( .fault(fault), .net(N466), .FEN(FEN[245]), .op(N466_t0) );
fim FAN_N466_1 ( .fault(fault), .net(N466), .FEN(FEN[246]), .op(N466_t1) );
fim FAN_N466_2 ( .fault(fault), .net(N466), .FEN(FEN[247]), .op(N466_t2) );
fim FAN_N466_3 ( .fault(fault), .net(N466), .FEN(FEN[248]), .op(N466_t3) );
fim FAN_N466_4 ( .fault(fault), .net(N466), .FEN(FEN[249]), .op(N466_t4) );
fim FAN_N466_5 ( .fault(fault), .net(N466), .FEN(FEN[250]), .op(N466_t5) );
fim FAN_N466_6 ( .fault(fault), .net(N466), .FEN(FEN[251]), .op(N466_t6) );
fim FAN_N466_7 ( .fault(fault), .net(N466), .FEN(FEN[252]), .op(N466_t7) );
fim FAN_N483_0 ( .fault(fault), .net(N483), .FEN(FEN[253]), .op(N483_t0) );
fim FAN_N483_1 ( .fault(fault), .net(N483), .FEN(FEN[254]), .op(N483_t1) );
fim FAN_N483_2 ( .fault(fault), .net(N483), .FEN(FEN[255]), .op(N483_t2) );
fim FAN_N483_3 ( .fault(fault), .net(N483), .FEN(FEN[256]), .op(N483_t3) );
fim FAN_N492_0 ( .fault(fault), .net(N492), .FEN(FEN[257]), .op(N492_t0) );
fim FAN_N492_1 ( .fault(fault), .net(N492), .FEN(FEN[258]), .op(N492_t1) );
fim FAN_N495_0 ( .fault(fault), .net(N495), .FEN(FEN[259]), .op(N495_t0) );
fim FAN_N495_1 ( .fault(fault), .net(N495), .FEN(FEN[260]), .op(N495_t1) );
fim FAN_N207_0 ( .fault(fault), .net(N207), .FEN(FEN[261]), .op(N207_t0) );
fim FAN_N207_1 ( .fault(fault), .net(N207), .FEN(FEN[262]), .op(N207_t1) );
fim FAN_N451_0 ( .fault(fault), .net(N451), .FEN(FEN[263]), .op(N451_t0) );
fim FAN_N451_1 ( .fault(fault), .net(N451), .FEN(FEN[264]), .op(N451_t1) );
fim FAN_N451_2 ( .fault(fault), .net(N451), .FEN(FEN[265]), .op(N451_t2) );
fim FAN_N451_3 ( .fault(fault), .net(N451), .FEN(FEN[266]), .op(N451_t3) );
fim FAN_N451_4 ( .fault(fault), .net(N451), .FEN(FEN[267]), .op(N451_t4) );
fim FAN_N451_5 ( .fault(fault), .net(N451), .FEN(FEN[268]), .op(N451_t5) );
fim FAN_N451_6 ( .fault(fault), .net(N451), .FEN(FEN[269]), .op(N451_t6) );
fim FAN_N451_7 ( .fault(fault), .net(N451), .FEN(FEN[270]), .op(N451_t7) );
fim FAN_N530_0 ( .fault(fault), .net(N530), .FEN(FEN[271]), .op(N530_t0) );
fim FAN_N530_1 ( .fault(fault), .net(N530), .FEN(FEN[272]), .op(N530_t1) );
fim FAN_N533_0 ( .fault(fault), .net(N533), .FEN(FEN[273]), .op(N533_t0) );
fim FAN_N533_1 ( .fault(fault), .net(N533), .FEN(FEN[274]), .op(N533_t1) );
fim FAN_N544_0 ( .fault(fault), .net(N544), .FEN(FEN[275]), .op(N544_t0) );
fim FAN_N544_1 ( .fault(fault), .net(N544), .FEN(FEN[276]), .op(N544_t1) );
fim FAN_N547_0 ( .fault(fault), .net(N547), .FEN(FEN[277]), .op(N547_t0) );
fim FAN_N547_1 ( .fault(fault), .net(N547), .FEN(FEN[278]), .op(N547_t1) );
fim FAN_N553_0 ( .fault(fault), .net(N553), .FEN(FEN[279]), .op(N553_t0) );
fim FAN_N553_1 ( .fault(fault), .net(N553), .FEN(FEN[280]), .op(N553_t1) );
fim FAN_N553_2 ( .fault(fault), .net(N553), .FEN(FEN[281]), .op(N553_t2) );
fim FAN_N246_0 ( .fault(fault), .net(N246), .FEN(FEN[282]), .op(N246_t0) );
fim FAN_N246_1 ( .fault(fault), .net(N246), .FEN(FEN[283]), .op(N246_t1) );
fim FAN_N246_2 ( .fault(fault), .net(N246), .FEN(FEN[284]), .op(N246_t2) );
fim FAN_N246_3 ( .fault(fault), .net(N246), .FEN(FEN[285]), .op(N246_t3) );
fim FAN_N246_4 ( .fault(fault), .net(N246), .FEN(FEN[286]), .op(N246_t4) );
fim FAN_N246_5 ( .fault(fault), .net(N246), .FEN(FEN[287]), .op(N246_t5) );
fim FAN_N246_6 ( .fault(fault), .net(N246), .FEN(FEN[288]), .op(N246_t6) );
fim FAN_N246_7 ( .fault(fault), .net(N246), .FEN(FEN[289]), .op(N246_t7) );
fim FAN_N557_0 ( .fault(fault), .net(N557), .FEN(FEN[290]), .op(N557_t0) );
fim FAN_N557_1 ( .fault(fault), .net(N557), .FEN(FEN[291]), .op(N557_t1) );
fim FAN_N557_2 ( .fault(fault), .net(N557), .FEN(FEN[292]), .op(N557_t2) );
fim FAN_N561_0 ( .fault(fault), .net(N561), .FEN(FEN[293]), .op(N561_t0) );
fim FAN_N561_1 ( .fault(fault), .net(N561), .FEN(FEN[294]), .op(N561_t1) );
fim FAN_N561_2 ( .fault(fault), .net(N561), .FEN(FEN[295]), .op(N561_t2) );
fim FAN_N565_0 ( .fault(fault), .net(N565), .FEN(FEN[296]), .op(N565_t0) );
fim FAN_N565_1 ( .fault(fault), .net(N565), .FEN(FEN[297]), .op(N565_t1) );
fim FAN_N565_2 ( .fault(fault), .net(N565), .FEN(FEN[298]), .op(N565_t2) );
fim FAN_N569_0 ( .fault(fault), .net(N569), .FEN(FEN[299]), .op(N569_t0) );
fim FAN_N569_1 ( .fault(fault), .net(N569), .FEN(FEN[300]), .op(N569_t1) );
fim FAN_N569_2 ( .fault(fault), .net(N569), .FEN(FEN[301]), .op(N569_t2) );
fim FAN_N573_0 ( .fault(fault), .net(N573), .FEN(FEN[302]), .op(N573_t0) );
fim FAN_N573_1 ( .fault(fault), .net(N573), .FEN(FEN[303]), .op(N573_t1) );
fim FAN_N573_2 ( .fault(fault), .net(N573), .FEN(FEN[304]), .op(N573_t2) );
fim FAN_N577_0 ( .fault(fault), .net(N577), .FEN(FEN[305]), .op(N577_t0) );
fim FAN_N577_1 ( .fault(fault), .net(N577), .FEN(FEN[306]), .op(N577_t1) );
fim FAN_N577_2 ( .fault(fault), .net(N577), .FEN(FEN[307]), .op(N577_t2) );
fim FAN_N581_0 ( .fault(fault), .net(N581), .FEN(FEN[308]), .op(N581_t0) );
fim FAN_N581_1 ( .fault(fault), .net(N581), .FEN(FEN[309]), .op(N581_t1) );
fim FAN_N581_2 ( .fault(fault), .net(N581), .FEN(FEN[310]), .op(N581_t2) );
fim FAN_N590_0 ( .fault(fault), .net(N590), .FEN(FEN[311]), .op(N590_t0) );
fim FAN_N590_1 ( .fault(fault), .net(N590), .FEN(FEN[312]), .op(N590_t1) );
fim FAN_N593_0 ( .fault(fault), .net(N593), .FEN(FEN[313]), .op(N593_t0) );
fim FAN_N593_1 ( .fault(fault), .net(N593), .FEN(FEN[314]), .op(N593_t1) );
fim FAN_N597_0 ( .fault(fault), .net(N597), .FEN(FEN[315]), .op(N597_t0) );
fim FAN_N597_1 ( .fault(fault), .net(N597), .FEN(FEN[316]), .op(N597_t1) );
fim FAN_N600_0 ( .fault(fault), .net(N600), .FEN(FEN[317]), .op(N600_t0) );
fim FAN_N600_1 ( .fault(fault), .net(N600), .FEN(FEN[318]), .op(N600_t1) );
fim FAN_N600_2 ( .fault(fault), .net(N600), .FEN(FEN[319]), .op(N600_t2) );
fim FAN_N600_3 ( .fault(fault), .net(N600), .FEN(FEN[320]), .op(N600_t3) );
fim FAN_N606_0 ( .fault(fault), .net(N606), .FEN(FEN[321]), .op(N606_t0) );
fim FAN_N606_1 ( .fault(fault), .net(N606), .FEN(FEN[322]), .op(N606_t1) );
fim FAN_N609_0 ( .fault(fault), .net(N609), .FEN(FEN[323]), .op(N609_t0) );
fim FAN_N609_1 ( .fault(fault), .net(N609), .FEN(FEN[324]), .op(N609_t1) );
fim FAN_N609_2 ( .fault(fault), .net(N609), .FEN(FEN[325]), .op(N609_t2) );
fim FAN_N609_3 ( .fault(fault), .net(N609), .FEN(FEN[326]), .op(N609_t3) );
fim FAN_N609_4 ( .fault(fault), .net(N609), .FEN(FEN[327]), .op(N609_t4) );
fim FAN_N616_0 ( .fault(fault), .net(N616), .FEN(FEN[328]), .op(N616_t0) );
fim FAN_N616_1 ( .fault(fault), .net(N616), .FEN(FEN[329]), .op(N616_t1) );
fim FAN_N619_0 ( .fault(fault), .net(N619), .FEN(FEN[330]), .op(N619_t0) );
fim FAN_N619_1 ( .fault(fault), .net(N619), .FEN(FEN[331]), .op(N619_t1) );
fim FAN_N619_2 ( .fault(fault), .net(N619), .FEN(FEN[332]), .op(N619_t2) );
fim FAN_N619_3 ( .fault(fault), .net(N619), .FEN(FEN[333]), .op(N619_t3) );
fim FAN_N625_0 ( .fault(fault), .net(N625), .FEN(FEN[334]), .op(N625_t0) );
fim FAN_N625_1 ( .fault(fault), .net(N625), .FEN(FEN[335]), .op(N625_t1) );
fim FAN_N628_0 ( .fault(fault), .net(N628), .FEN(FEN[336]), .op(N628_t0) );
fim FAN_N628_1 ( .fault(fault), .net(N628), .FEN(FEN[337]), .op(N628_t1) );
fim FAN_N632_0 ( .fault(fault), .net(N632), .FEN(FEN[338]), .op(N632_t0) );
fim FAN_N632_1 ( .fault(fault), .net(N632), .FEN(FEN[339]), .op(N632_t1) );
fim FAN_N635_0 ( .fault(fault), .net(N635), .FEN(FEN[340]), .op(N635_t0) );
fim FAN_N635_1 ( .fault(fault), .net(N635), .FEN(FEN[341]), .op(N635_t1) );
fim FAN_N635_2 ( .fault(fault), .net(N635), .FEN(FEN[342]), .op(N635_t2) );
fim FAN_N635_3 ( .fault(fault), .net(N635), .FEN(FEN[343]), .op(N635_t3) );
fim FAN_N641_0 ( .fault(fault), .net(N641), .FEN(FEN[344]), .op(N641_t0) );
fim FAN_N641_1 ( .fault(fault), .net(N641), .FEN(FEN[345]), .op(N641_t1) );
fim FAN_N644_0 ( .fault(fault), .net(N644), .FEN(FEN[346]), .op(N644_t0) );
fim FAN_N644_1 ( .fault(fault), .net(N644), .FEN(FEN[347]), .op(N644_t1) );
fim FAN_N644_2 ( .fault(fault), .net(N644), .FEN(FEN[348]), .op(N644_t2) );
fim FAN_N644_3 ( .fault(fault), .net(N644), .FEN(FEN[349]), .op(N644_t3) );
fim FAN_N644_4 ( .fault(fault), .net(N644), .FEN(FEN[350]), .op(N644_t4) );
fim FAN_N651_0 ( .fault(fault), .net(N651), .FEN(FEN[351]), .op(N651_t0) );
fim FAN_N651_1 ( .fault(fault), .net(N651), .FEN(FEN[352]), .op(N651_t1) );
fim FAN_N654_0 ( .fault(fault), .net(N654), .FEN(FEN[353]), .op(N654_t0) );
fim FAN_N654_1 ( .fault(fault), .net(N654), .FEN(FEN[354]), .op(N654_t1) );
fim FAN_N654_2 ( .fault(fault), .net(N654), .FEN(FEN[355]), .op(N654_t2) );
fim FAN_N654_3 ( .fault(fault), .net(N654), .FEN(FEN[356]), .op(N654_t3) );
fim FAN_N261_0 ( .fault(fault), .net(N261), .FEN(FEN[357]), .op(N261_t0) );
fim FAN_N261_1 ( .fault(fault), .net(N261), .FEN(FEN[358]), .op(N261_t1) );
fim FAN_N261_2 ( .fault(fault), .net(N261), .FEN(FEN[359]), .op(N261_t2) );
fim FAN_N261_3 ( .fault(fault), .net(N261), .FEN(FEN[360]), .op(N261_t3) );
fim FAN_N261_4 ( .fault(fault), .net(N261), .FEN(FEN[361]), .op(N261_t4) );
fim FAN_N662_0 ( .fault(fault), .net(N662), .FEN(FEN[362]), .op(N662_t0) );
fim FAN_N662_1 ( .fault(fault), .net(N662), .FEN(FEN[363]), .op(N662_t1) );
fim FAN_N228_0 ( .fault(fault), .net(N228), .FEN(FEN[364]), .op(N228_t0) );
fim FAN_N228_1 ( .fault(fault), .net(N228), .FEN(FEN[365]), .op(N228_t1) );
fim FAN_N228_2 ( .fault(fault), .net(N228), .FEN(FEN[366]), .op(N228_t2) );
fim FAN_N228_3 ( .fault(fault), .net(N228), .FEN(FEN[367]), .op(N228_t3) );
fim FAN_N228_4 ( .fault(fault), .net(N228), .FEN(FEN[368]), .op(N228_t4) );
fim FAN_N228_5 ( .fault(fault), .net(N228), .FEN(FEN[369]), .op(N228_t5) );
fim FAN_N228_6 ( .fault(fault), .net(N228), .FEN(FEN[370]), .op(N228_t6) );
fim FAN_N228_7 ( .fault(fault), .net(N228), .FEN(FEN[371]), .op(N228_t7) );
fim FAN_N665_0 ( .fault(fault), .net(N665), .FEN(FEN[372]), .op(N665_t0) );
fim FAN_N665_1 ( .fault(fault), .net(N665), .FEN(FEN[373]), .op(N665_t1) );
fim FAN_N665_2 ( .fault(fault), .net(N665), .FEN(FEN[374]), .op(N665_t2) );
fim FAN_N237_0 ( .fault(fault), .net(N237), .FEN(FEN[375]), .op(N237_t0) );
fim FAN_N237_1 ( .fault(fault), .net(N237), .FEN(FEN[376]), .op(N237_t1) );
fim FAN_N237_2 ( .fault(fault), .net(N237), .FEN(FEN[377]), .op(N237_t2) );
fim FAN_N237_3 ( .fault(fault), .net(N237), .FEN(FEN[378]), .op(N237_t3) );
fim FAN_N237_4 ( .fault(fault), .net(N237), .FEN(FEN[379]), .op(N237_t4) );
fim FAN_N237_5 ( .fault(fault), .net(N237), .FEN(FEN[380]), .op(N237_t5) );
fim FAN_N237_6 ( .fault(fault), .net(N237), .FEN(FEN[381]), .op(N237_t6) );
fim FAN_N237_7 ( .fault(fault), .net(N237), .FEN(FEN[382]), .op(N237_t7) );
fim FAN_N670_0 ( .fault(fault), .net(N670), .FEN(FEN[383]), .op(N670_t0) );
fim FAN_N670_1 ( .fault(fault), .net(N670), .FEN(FEN[384]), .op(N670_t1) );
fim FAN_N673_0 ( .fault(fault), .net(N673), .FEN(FEN[385]), .op(N673_t0) );
fim FAN_N673_1 ( .fault(fault), .net(N673), .FEN(FEN[386]), .op(N673_t1) );
fim FAN_N673_2 ( .fault(fault), .net(N673), .FEN(FEN[387]), .op(N673_t2) );
fim FAN_N678_0 ( .fault(fault), .net(N678), .FEN(FEN[388]), .op(N678_t0) );
fim FAN_N678_1 ( .fault(fault), .net(N678), .FEN(FEN[389]), .op(N678_t1) );
fim FAN_N678_2 ( .fault(fault), .net(N678), .FEN(FEN[390]), .op(N678_t2) );
fim FAN_N682_0 ( .fault(fault), .net(N682), .FEN(FEN[391]), .op(N682_t0) );
fim FAN_N682_1 ( .fault(fault), .net(N682), .FEN(FEN[392]), .op(N682_t1) );
fim FAN_N682_2 ( .fault(fault), .net(N682), .FEN(FEN[393]), .op(N682_t2) );
fim FAN_N687_0 ( .fault(fault), .net(N687), .FEN(FEN[394]), .op(N687_t0) );
fim FAN_N687_1 ( .fault(fault), .net(N687), .FEN(FEN[395]), .op(N687_t1) );
fim FAN_N687_2 ( .fault(fault), .net(N687), .FEN(FEN[396]), .op(N687_t2) );
fim FAN_N687_3 ( .fault(fault), .net(N687), .FEN(FEN[397]), .op(N687_t3) );
fim FAN_N692_0 ( .fault(fault), .net(N692), .FEN(FEN[398]), .op(N692_t0) );
fim FAN_N692_1 ( .fault(fault), .net(N692), .FEN(FEN[399]), .op(N692_t1) );
fim FAN_N692_2 ( .fault(fault), .net(N692), .FEN(FEN[400]), .op(N692_t2) );
fim FAN_N697_0 ( .fault(fault), .net(N697), .FEN(FEN[401]), .op(N697_t0) );
fim FAN_N697_1 ( .fault(fault), .net(N697), .FEN(FEN[402]), .op(N697_t1) );
fim FAN_N700_0 ( .fault(fault), .net(N700), .FEN(FEN[403]), .op(N700_t0) );
fim FAN_N700_1 ( .fault(fault), .net(N700), .FEN(FEN[404]), .op(N700_t1) );
fim FAN_N700_2 ( .fault(fault), .net(N700), .FEN(FEN[405]), .op(N700_t2) );
fim FAN_N705_0 ( .fault(fault), .net(N705), .FEN(FEN[406]), .op(N705_t0) );
fim FAN_N705_1 ( .fault(fault), .net(N705), .FEN(FEN[407]), .op(N705_t1) );
fim FAN_N708_0 ( .fault(fault), .net(N708), .FEN(FEN[408]), .op(N708_t0) );
fim FAN_N708_1 ( .fault(fault), .net(N708), .FEN(FEN[409]), .op(N708_t1) );
fim FAN_N708_2 ( .fault(fault), .net(N708), .FEN(FEN[410]), .op(N708_t2) );
fim FAN_N713_0 ( .fault(fault), .net(N713), .FEN(FEN[411]), .op(N713_t0) );
fim FAN_N713_1 ( .fault(fault), .net(N713), .FEN(FEN[412]), .op(N713_t1) );
fim FAN_N713_2 ( .fault(fault), .net(N713), .FEN(FEN[413]), .op(N713_t2) );
fim FAN_N717_0 ( .fault(fault), .net(N717), .FEN(FEN[414]), .op(N717_t0) );
fim FAN_N717_1 ( .fault(fault), .net(N717), .FEN(FEN[415]), .op(N717_t1) );
fim FAN_N717_2 ( .fault(fault), .net(N717), .FEN(FEN[416]), .op(N717_t2) );
fim FAN_N722_0 ( .fault(fault), .net(N722), .FEN(FEN[417]), .op(N722_t0) );
fim FAN_N722_1 ( .fault(fault), .net(N722), .FEN(FEN[418]), .op(N722_t1) );
fim FAN_N722_2 ( .fault(fault), .net(N722), .FEN(FEN[419]), .op(N722_t2) );
fim FAN_N722_3 ( .fault(fault), .net(N722), .FEN(FEN[420]), .op(N722_t3) );
fim FAN_N727_0 ( .fault(fault), .net(N727), .FEN(FEN[421]), .op(N727_t0) );
fim FAN_N727_1 ( .fault(fault), .net(N727), .FEN(FEN[422]), .op(N727_t1) );
fim FAN_N727_2 ( .fault(fault), .net(N727), .FEN(FEN[423]), .op(N727_t2) );
fim FAN_N773_0 ( .fault(fault), .net(N773), .FEN(FEN[424]), .op(N773_t0) );
fim FAN_N773_1 ( .fault(fault), .net(N773), .FEN(FEN[425]), .op(N773_t1) );
fim FAN_N773_2 ( .fault(fault), .net(N773), .FEN(FEN[426]), .op(N773_t2) );
fim FAN_N778_0 ( .fault(fault), .net(N778), .FEN(FEN[427]), .op(N778_t0) );
fim FAN_N778_1 ( .fault(fault), .net(N778), .FEN(FEN[428]), .op(N778_t1) );
fim FAN_N782_0 ( .fault(fault), .net(N782), .FEN(FEN[429]), .op(N782_t0) );
fim FAN_N782_1 ( .fault(fault), .net(N782), .FEN(FEN[430]), .op(N782_t1) );
fim FAN_N219_0 ( .fault(fault), .net(N219), .FEN(FEN[431]), .op(N219_t0) );
fim FAN_N219_1 ( .fault(fault), .net(N219), .FEN(FEN[432]), .op(N219_t1) );
fim FAN_N219_2 ( .fault(fault), .net(N219), .FEN(FEN[433]), .op(N219_t2) );
fim FAN_N219_3 ( .fault(fault), .net(N219), .FEN(FEN[434]), .op(N219_t3) );
fim FAN_N219_4 ( .fault(fault), .net(N219), .FEN(FEN[435]), .op(N219_t4) );
fim FAN_N219_5 ( .fault(fault), .net(N219), .FEN(FEN[436]), .op(N219_t5) );
fim FAN_N219_6 ( .fault(fault), .net(N219), .FEN(FEN[437]), .op(N219_t6) );
fim FAN_N219_7 ( .fault(fault), .net(N219), .FEN(FEN[438]), .op(N219_t7) );
fim FAN_N796_0 ( .fault(fault), .net(N796), .FEN(FEN[439]), .op(N796_t0) );
fim FAN_N796_1 ( .fault(fault), .net(N796), .FEN(FEN[440]), .op(N796_t1) );
fim FAN_N796_2 ( .fault(fault), .net(N796), .FEN(FEN[441]), .op(N796_t2) );
fim FAN_N796_3 ( .fault(fault), .net(N796), .FEN(FEN[442]), .op(N796_t3) );
fim FAN_N796_4 ( .fault(fault), .net(N796), .FEN(FEN[443]), .op(N796_t4) );
fim FAN_N815_0 ( .fault(fault), .net(N815), .FEN(FEN[444]), .op(N815_t0) );
fim FAN_N815_1 ( .fault(fault), .net(N815), .FEN(FEN[445]), .op(N815_t1) );
fim FAN_N815_2 ( .fault(fault), .net(N815), .FEN(FEN[446]), .op(N815_t2) );
fim FAN_N819_0 ( .fault(fault), .net(N819), .FEN(FEN[447]), .op(N819_t0) );
fim FAN_N819_1 ( .fault(fault), .net(N819), .FEN(FEN[448]), .op(N819_t1) );
fim FAN_N822_0 ( .fault(fault), .net(N822), .FEN(FEN[449]), .op(N822_t0) );
fim FAN_N822_1 ( .fault(fault), .net(N822), .FEN(FEN[450]), .op(N822_t1) );
initial begin
    FEN <= {450'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {450'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,450'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,450'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN <= {FEN[449:0], FEN[450]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
// EndFaultModel

//Anchor
nand NAND4_1 (N269, N1_t0, N8_t0, N13_t0, N17_t0);
nand NAND4_2 (N270, N1_t1, N26_t0, N13_t1, N17_t1);
and AND3_3 (N273, N29_t0, N36_t0, N42_t0);
and AND3_4 (N276, N1_t2, N26_t1, N51_t0);
nand NAND4_5 (N279, N1_t3, N8_t1, N51_t1, N17_t2);
nand NAND4_6 (N280, N1_t4, N8_t2, N13_t2, N55_t0);
nand NAND4_7 (N284, N59_t0, N42_t1, N68_t0, N72_t);
nand NAND2_8 (N285, N29_t1, N68_t1);
nand NAND3_9 (N286, N59_t1, N68_t2, N74_t);
and AND3_10 (N287, N29_t2, N75_t0, N80_t0);
and AND3_11 (N290, N29_t3, N75_t1, N42_t2);
and AND3_12 (N291, N29_t4, N36_t1, N80_t1);
and AND3_13 (N292, N29_t5, N36_t2, N42_t3);
and AND3_14 (N293, N59_t2, N75_t2, N80_t2);
and AND3_15 (N294, N59_t3, N75_t3, N42_t4);
and AND3_16 (N295, N59_t4, N36_t3, N80_t3);
and AND3_17 (N296, N59_t5, N36_t4, N42_t5);
and AND2_18 (N297, N85_t, N86_t);
or OR2_19 (N298, N87_t, N88_t);
nand NAND2_20 (N301, N91_t0, N96_t0);
or OR2_21 (N302, N91_t1, N96_t1);
nand NAND2_22 (N303, N101_t0, N106_t0);
or OR2_23 (N304, N101_t1, N106_t1);
nand NAND2_24 (N305, N111_t0, N116_t0);
or OR2_25 (N306, N111_t1, N116_t1);
nand NAND2_26 (N307, N121_t0, N126_t0);
or OR2_27 (N308, N121_t1, N126_t1);
and AND2_28 (N309, N8_t3, N138_t0);
not NOT1_29 (N310, N268_t);
and AND2_30 (N316, N51_t2, N138_t1);
and AND2_31 (N317, N17_t3, N138_t2);
and AND2_32 (N318, N152_t, N138_t3);
nand NAND2_33 (N319, N59_t6, N156_t0);
nor NOR2_34 (N322, N17_t4, N42_t6);
and AND2_35 (N323, N17_t5, N42_t7);
nand NAND2_36 (N324, N159_t0, N165_t0);
or OR2_37 (N325, N159_t1, N165_t1);
nand NAND2_38 (N326, N171_t0, N177_t0);
or OR2_39 (N327, N171_t1, N177_t1);
nand NAND2_40 (N328, N183_t0, N189_t0);
or OR2_41 (N329, N183_t1, N189_t1);
nand NAND2_42 (N330, N195_t0, N201_t0);
or OR2_43 (N331, N195_t1, N201_t1);
and AND2_44 (N332, N210_t0, N91_t2);
and AND2_45 (N333, N210_t1, N96_t2);
and AND2_46 (N334, N210_t2, N101_t2);
and AND2_47 (N335, N210_t3, N106_t2);
and AND2_48 (N336, N210_t4, N111_t2);
and AND2_49 (N337, N255_t0, N259_t);
and AND2_50 (N338, N210_t5, N116_t2);
and AND2_51 (N339, N255_t1, N260_t);
and AND2_52 (N340, N210_t6, N121_t2);
and AND2_53 (N341, N255_t2, N267_t);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273_t0);
or OR2_56 (N344, N270_t0, N273_t1);
not NOT1_57 (N345, N276_t0);
not NOT1_58 (N346, N276_t1);
not NOT1_59 (N347, N279);
nor NOR2_60 (N348, N280_t0, N284);
or OR2_61 (N349, N280_t1, N285);
or OR2_62 (N350, N280_t2, N286);
not NOT1_63 (N351, N293);
not NOT1_64 (N352, N294);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89_t, N298_t0);
and AND2_68 (N356, N90_t, N298_t1);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
not NOT1_73 (N369, N310_t0);
nor NOR2_74 (N375, N322, N323);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270_t1, N343);
not NOT1_84 (N393, N345);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73_t);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357_t0);
not NOT1_91 (N405, N360_t0);
and AND2_92 (N406, N357_t1, N360_t1);
not NOT1_93 (N407, N363_t0);
not NOT1_94 (N408, N366_t0);
and AND2_95 (N409, N363_t1, N366_t1);
nand NAND2_96 (N410, N347, N352);
not NOT1_97 (N411, N376_t0);
not NOT1_98 (N412, N379_t0);
and AND2_99 (N413, N376_t1, N379_t1);
not NOT1_100 (N414, N382_t0);
not NOT1_101 (N415, N385_t0);
and AND2_102 (N416, N382_t1, N385_t1);
and AND2_103 (N417, N210_t7, N369_t0);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
and AND3_113 (N427, N319_t0, N393_t0, N55_t1);
and AND3_114 (N432, N393_t1, N17_t6, N287_t0);
nand NAND3_115 (N437, N393_t2, N287_t1, N55_t2);
nand NAND4_116 (N442, N375, N59_t7, N156_t1, N393_t3);
nand NAND3_117 (N443, N393_t4, N319_t1, N17_t7);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
nand NAND2_128 (N466, N442, N410);
and AND2_129 (N475, N143_t0, N427_t0);
and AND2_130 (N476, N310_t1, N432_t0);
and AND2_131 (N477, N146_t0, N427_t1);
and AND2_132 (N478, N310_t2, N432_t1);
and AND2_133 (N479, N149_t0, N427_t2);
and AND2_134 (N480, N310_t3, N432_t2);
and AND2_135 (N481, N153_t0, N427_t3);
and AND2_136 (N482, N310_t4, N432_t3);
nand NAND2_137 (N483, N443, N1_t5);
or OR2_138 (N488, N369_t1, N437_t0);
or OR2_139 (N489, N369_t2, N437_t1);
or OR2_140 (N490, N369_t3, N437_t2);
or OR2_141 (N491, N369_t4, N437_t3);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130_t0, N460_t0);
or OR2_145 (N499, N130_t1, N460_t1);
nand NAND2_146 (N500, N463_t0, N135_t0);
or OR2_147 (N501, N463_t1, N135_t1);
and AND2_148 (N502, N91_t3, N466_t0);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96_t3, N466_t1);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101_t3, N466_t2);
nor NOR2_153 (N507, N479, N480);
and AND2_154 (N508, N106_t3, N466_t3);
nor NOR2_155 (N509, N481, N482);
and AND2_156 (N510, N143_t1, N483_t0);
and AND2_157 (N511, N111_t3, N466_t4);
and AND2_158 (N512, N146_t1, N483_t1);
and AND2_159 (N513, N116_t3, N466_t5);
and AND2_160 (N514, N149_t1, N483_t2);
and AND2_161 (N515, N121_t3, N466_t6);
and AND2_162 (N516, N153_t1, N483_t3);
and AND2_163 (N517, N126_t2, N466_t7);
nand NAND2_164 (N518, N130_t2, N492_t0);
or OR2_165 (N519, N130_t3, N492_t1);
nand NAND2_166 (N520, N495_t0, N207_t0);
or OR2_167 (N521, N495_t1, N207_t1);
and AND2_168 (N522, N451_t0, N159_t2);
and AND2_169 (N523, N451_t1, N165_t2);
and AND2_170 (N524, N451_t2, N171_t2);
and AND2_171 (N525, N451_t3, N177_t2);
and AND2_172 (N526, N451_t4, N183_t2);
nand NAND2_173 (N527, N451_t5, N189_t2);
nand NAND2_174 (N528, N451_t6, N195_t2);
nand NAND2_175 (N529, N451_t7, N201_t2);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
nor NOR2_182 (N540, N510, N511);
nor NOR2_183 (N541, N512, N513);
nor NOR2_184 (N542, N514, N515);
nor NOR2_185 (N543, N516, N517);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530_t0);
not NOT1_189 (N551, N533_t0);
and AND2_190 (N552, N530_t1, N533_t1);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
nand NAND2_193 (N561, N538, N507);
nand NAND2_194 (N565, N539, N509);
nand NAND2_195 (N569, N488, N540);
nand NAND2_196 (N573, N489, N541);
nand NAND2_197 (N577, N490, N542);
nand NAND2_198 (N581, N491, N543);
not NOT1_199 (N585, N544_t0);
not NOT1_200 (N586, N547_t0);
and AND2_201 (N587, N544_t1, N547_t1);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
nand NAND2_204 (N590, N553_t0, N159_t3);
or OR2_205 (N593, N553_t1, N159_t4);
and AND2_206 (N596, N246_t0, N553_t2);
nand NAND2_207 (N597, N557_t0, N165_t3);
or OR2_208 (N600, N557_t1, N165_t4);
and AND2_209 (N605, N246_t1, N557_t2);
nand NAND2_210 (N606, N561_t0, N171_t3);
or OR2_211 (N609, N561_t1, N171_t4);
and AND2_212 (N615, N246_t2, N561_t2);
nand NAND2_213 (N616, N565_t0, N177_t3);
or OR2_214 (N619, N565_t1, N177_t4);
and AND2_215 (N624, N246_t3, N565_t2);
nand NAND2_216 (N625, N569_t0, N183_t3);
or OR2_217 (N628, N569_t1, N183_t4);
and AND2_218 (N631, N246_t4, N569_t2);
nand NAND2_219 (N632, N573_t0, N189_t3);
or OR2_220 (N635, N573_t1, N189_t4);
and AND2_221 (N640, N246_t5, N573_t2);
nand NAND2_222 (N641, N577_t0, N195_t3);
or OR2_223 (N644, N577_t1, N195_t4);
and AND2_224 (N650, N246_t6, N577_t2);
nand NAND2_225 (N651, N581_t0, N201_t3);
or OR2_226 (N654, N581_t1, N201_t4);
and AND2_227 (N659, N246_t7, N581_t2);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590_t0);
and AND2_231 (N665, N593_t0, N590_t1);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597_t0);
and AND2_234 (N673, N600_t0, N597_t1);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606_t0);
and AND2_237 (N682, N609_t0, N606_t1);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616_t0);
and AND2_240 (N692, N619_t0, N616_t1);
nor NOR2_241 (N696, N624, N525);
not NOT1_242 (N697, N625_t0);
and AND2_243 (N700, N628_t0, N625_t1);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632_t0);
and AND2_246 (N708, N635_t0, N632_t1);
nor NOR2_247 (N712, N337, N640);
not NOT1_248 (N713, N641_t0);
and AND2_249 (N717, N644_t0, N641_t1);
nor NOR2_250 (N721, N339, N650);
not NOT1_251 (N722, N651_t0);
and AND2_252 (N727, N654_t0, N651_t1);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654_t1, N261_t0);
nand NAND3_255 (N733, N644_t1, N654_t2, N261_t1);
nand NAND4_256 (N734, N635_t1, N644_t2, N654_t3, N261_t2);
not NOT1_257 (N735, N662_t0);
and AND2_258 (N736, N228_t0, N665_t0);
and AND2_259 (N737, N237_t0, N662_t1);
not NOT1_260 (N738, N670_t0);
and AND2_261 (N739, N228_t1, N673_t0);
and AND2_262 (N740, N237_t1, N670_t1);
not NOT1_263 (N741, N678_t0);
and AND2_264 (N742, N228_t2, N682_t0);
and AND2_265 (N743, N237_t2, N678_t1);
not NOT1_266 (N744, N687_t0);
and AND2_267 (N745, N228_t3, N692_t0);
and AND2_268 (N746, N237_t3, N687_t1);
not NOT1_269 (N747, N697_t0);
and AND2_270 (N748, N228_t4, N700_t0);
and AND2_271 (N749, N237_t4, N697_t1);
not NOT1_272 (N750, N705_t0);
and AND2_273 (N751, N228_t5, N708_t0);
and AND2_274 (N752, N237_t5, N705_t1);
not NOT1_275 (N753, N713_t0);
and AND2_276 (N754, N228_t6, N717_t0);
and AND2_277 (N755, N237_t6, N713_t1);
not NOT1_278 (N756, N722_t0);
nor NOR2_279 (N757, N727_t0, N261_t3);
and AND2_280 (N758, N727_t1, N261_t4);
and AND2_281 (N759, N228_t7, N727_t2);
and AND2_282 (N760, N237_t7, N722_t1);
nand NAND2_283 (N761, N644_t3, N722_t2);
nand NAND2_284 (N762, N635_t2, N713_t2);
nand NAND3_285 (N763, N635_t3, N644_t4, N722_t3);
nand NAND2_286 (N764, N609_t1, N687_t2);
nand NAND2_287 (N765, N600_t1, N678_t2);
nand NAND3_288 (N766, N600_t2, N609_t2, N687_t3);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
nand NAND4_295 (N773, N750, N762, N763, N734);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
nor NOR2_303 (N788, N700_t1, N773_t0);
and AND2_304 (N789, N700_t2, N773_t1);
nor NOR2_305 (N790, N708_t1, N778_t0);
and AND2_306 (N791, N708_t2, N778_t1);
nor NOR2_307 (N792, N717_t1, N782_t0);
and AND2_308 (N793, N717_t2, N782_t1);
and AND2_309 (N794, N219_t0, N786);
nand NAND2_310 (N795, N628_t1, N773_t2);
nand NAND2_311 (N796, N795, N747);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
nor NOR2_316 (N806, N692_t1, N796_t0);
and AND2_317 (N807, N692_t2, N796_t1);
and AND2_318 (N808, N219_t1, N802);
and AND2_319 (N809, N219_t2, N803);
and AND2_320 (N810, N219_t3, N804);
nand NAND4_321 (N811, N805, N787, N731, N529);
nand NAND2_322 (N812, N619_t1, N796_t2);
nand NAND3_323 (N813, N609_t3, N619_t2, N796_t3);
nand NAND4_324 (N814, N600_t3, N609_t4, N619_t3, N796_t4);
nand NAND4_325 (N815, N738, N765, N766, N814);
nand NAND3_326 (N819, N741, N764, N813);
nand NAND2_327 (N822, N744, N812);
nor NOR2_328 (N825, N806, N807);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
nor NOR2_333 (N830, N665_t1, N815_t0);
and AND2_334 (N831, N665_t2, N815_t1);
nor NOR2_335 (N832, N673_t1, N819_t0);
and AND2_336 (N833, N673_t2, N819_t1);
nor NOR2_337 (N834, N682_t1, N822_t0);
and AND2_338 (N835, N682_t2, N822_t1);
and AND2_339 (N836, N219_t4, N825);
nand NAND3_340 (N837, N826, N777, N704);
nand NAND4_341 (N838, N827, N781, N712, N527);
nand NAND4_342 (N839, N828, N785, N721, N528);
not NOT1_343 (N840, N829);
nand NAND2_344 (N841, N815_t2, N593_t1);
nor NOR2_345 (N842, N830, N831);
nor NOR2_346 (N843, N832, N833);
nor NOR2_347 (N844, N834, N835);
nor NOR2_348 (N845, N334, N836);
not NOT1_349 (N846, N837);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
and AND2_352 (N849, N735, N841);
buf BUFF1_353 (N850, N840);
and AND2_354 (N851, N219_t5, N842);
and AND2_355 (N852, N219_t6, N843);
and AND2_356 (N853, N219_t7, N844);
nand NAND3_357 (N854, N845, N772, N696);
not NOT1_358 (N855, N846);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
not NOT1_361 (N858, N849);
nor NOR2_362 (N859, N417, N851);
nor NOR2_363 (N860, N332, N852);
nor NOR2_364 (N861, N333, N853);
not NOT1_365 (N862, N854);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
nand NAND3_370 (N867, N859, N769, N669);
nand NAND3_371 (N868, N860, N770, N677);
nand NAND3_372 (N869, N861, N771, N686);
not NOT1_373 (N870, N862);
not NOT1_374 (N871, N867);
not NOT1_375 (N872, N868);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
not NOT1_378 (N875, N871);
not NOT1_379 (N876, N872);
not NOT1_380 (N877, N873);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

endmodule
