/* 
    BIST Controller

    Wraps together all the blocks of BIST functionality
*/

module bist_c(
);
    
endmodule