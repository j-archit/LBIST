/* 
    Test Pattern Generator

    Consists of 
    1.

*/

module tpg
(
);
    
endmodule