// Verilog
// c6288
// Ninputs 32
// Noutputs 32
// NtotalGates 2416
// AND2 256
// NOT1 32
// NOR2 2128

module c6288f (INC,END,clk,rst,N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,
              N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,
              N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,
              N511,N528,N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,
              N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,
              N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,
              N6270,N6280,N6287,N6288);

input N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,
      N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,
      N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,
      N511,N528;

output N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,
       N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,
       N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,
       N6287,N6288;

wire N546,N549,N552,N555,N558,N561,N564,N567,N570,N573,
     N576,N579,N582,N585,N588,N591,N594,N597,N600,N603,
     N606,N609,N612,N615,N618,N621,N624,N627,N630,N633,
     N636,N639,N642,N645,N648,N651,N654,N657,N660,N663,
     N666,N669,N672,N675,N678,N681,N684,N687,N690,N693,
     N696,N699,N702,N705,N708,N711,N714,N717,N720,N723,
     N726,N729,N732,N735,N738,N741,N744,N747,N750,N753,
     N756,N759,N762,N765,N768,N771,N774,N777,N780,N783,
     N786,N789,N792,N795,N798,N801,N804,N807,N810,N813,
     N816,N819,N822,N825,N828,N831,N834,N837,N840,N843,
     N846,N849,N852,N855,N858,N861,N864,N867,N870,N873,
     N876,N879,N882,N885,N888,N891,N894,N897,N900,N903,
     N906,N909,N912,N915,N918,N921,N924,N927,N930,N933,
     N936,N939,N942,N945,N948,N951,N954,N957,N960,N963,
     N966,N969,N972,N975,N978,N981,N984,N987,N990,N993,
     N996,N999,N1002,N1005,N1008,N1011,N1014,N1017,N1020,N1023,
     N1026,N1029,N1032,N1035,N1038,N1041,N1044,N1047,N1050,N1053,
     N1056,N1059,N1062,N1065,N1068,N1071,N1074,N1077,N1080,N1083,
     N1086,N1089,N1092,N1095,N1098,N1101,N1104,N1107,N1110,N1113,
     N1116,N1119,N1122,N1125,N1128,N1131,N1134,N1137,N1140,N1143,
     N1146,N1149,N1152,N1155,N1158,N1161,N1164,N1167,N1170,N1173,
     N1176,N1179,N1182,N1185,N1188,N1191,N1194,N1197,N1200,N1203,
     N1206,N1209,N1212,N1215,N1218,N1221,N1224,N1227,N1230,N1233,
     N1236,N1239,N1242,N1245,N1248,N1251,N1254,N1257,N1260,N1263,
     N1266,N1269,N1272,N1275,N1278,N1281,N1284,N1287,N1290,N1293,
     N1296,N1299,N1302,N1305,N1308,N1311,N1315,N1319,N1323,N1327,
     N1331,N1335,N1339,N1343,N1347,N1351,N1355,N1359,N1363,N1367,
     N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,
     N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,
     N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,
     N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,N1425,N1428,
     N1431,N1434,N1437,N1440,N1443,N1446,N1450,N1454,N1458,N1462,
     N1466,N1470,N1474,N1478,N1482,N1486,N1490,N1494,N1498,N1502,
     N1506,N1507,N1508,N1511,N1512,N1513,N1516,N1517,N1518,N1521,
     N1522,N1523,N1526,N1527,N1528,N1531,N1532,N1533,N1536,N1537,
     N1538,N1541,N1542,N1543,N1546,N1547,N1548,N1551,N1552,N1553,
     N1556,N1557,N1558,N1561,N1562,N1563,N1566,N1567,N1568,N1571,
     N1572,N1573,N1576,N1577,N1578,N1582,N1585,N1588,N1591,N1594,
     N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,N1621,N1624,
     N1628,N1632,N1636,N1640,N1644,N1648,N1652,N1656,N1660,N1664,
     N1668,N1672,N1676,N1680,N1684,N1685,N1686,N1687,N1688,N1689,
     N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,
     N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,
     N1710,N1711,N1712,N1713,N1714,N1717,N1720,N1723,N1726,N1729,
     N1732,N1735,N1738,N1741,N1744,N1747,N1750,N1753,N1756,N1759,
     N1763,N1767,N1771,N1775,N1779,N1783,N1787,N1791,N1795,N1799,
     N1803,N1807,N1811,N1815,N1819,N1820,N1821,N1824,N1825,N1826,
     N1829,N1830,N1831,N1834,N1835,N1836,N1839,N1840,N1841,N1844,
     N1845,N1846,N1849,N1850,N1851,N1854,N1855,N1856,N1859,N1860,
     N1861,N1864,N1865,N1866,N1869,N1870,N1871,N1874,N1875,N1876,
     N1879,N1880,N1881,N1884,N1885,N1886,N1889,N1890,N1891,N1894,
     N1897,N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,
     N1929,N1932,N1935,N1938,N1941,N1945,N1946,N1947,N1951,N1955,
     N1959,N1963,N1967,N1971,N1975,N1979,N1983,N1987,N1991,N1995,
     N1999,N2000,N2001,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
     N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,
     N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,
     N2033,N2037,N2040,N2043,N2046,N2049,N2052,N2055,N2058,N2061,
     N2064,N2067,N2070,N2073,N2076,N2080,N2081,N2082,N2085,N2089,
     N2093,N2097,N2101,N2105,N2109,N2113,N2117,N2121,N2125,N2129,
     N2133,N2137,N2138,N2139,N2142,N2145,N2149,N2150,N2151,N2154,
     N2155,N2156,N2159,N2160,N2161,N2164,N2165,N2166,N2169,N2170,
     N2171,N2174,N2175,N2176,N2179,N2180,N2181,N2184,N2185,N2186,
     N2189,N2190,N2191,N2194,N2195,N2196,N2199,N2200,N2201,N2204,
     N2205,N2206,N2209,N2210,N2211,N2214,N2217,N2221,N2222,N2224,
     N2227,N2230,N2233,N2236,N2239,N2242,N2245,N2248,N2251,N2254,
     N2257,N2260,N2264,N2265,N2266,N2269,N2273,N2277,N2281,N2285,
     N2289,N2293,N2297,N2301,N2305,N2309,N2313,N2317,N2318,N2319,
     N2322,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,
     N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
     N2345,N2346,N2347,N2348,N2349,N2350,N2353,N2357,N2358,N2359,
     N2362,N2365,N2368,N2371,N2374,N2377,N2380,N2383,N2386,N2389,
     N2392,N2395,N2398,N2402,N2403,N2404,N2407,N2410,N2414,N2418,
     N2422,N2426,N2430,N2434,N2438,N2442,N2446,N2450,N2454,N2458,
     N2462,N2463,N2464,N2467,N2470,N2474,N2475,N2476,N2477,N2478,
     N2481,N2482,N2483,N2486,N2487,N2488,N2491,N2492,N2493,N2496,
     N2497,N2498,N2501,N2502,N2503,N2506,N2507,N2508,N2511,N2512,
     N2513,N2516,N2517,N2518,N2521,N2522,N2523,N2526,N2527,N2528,
     N2531,N2532,N2533,N2536,N2539,N2543,N2544,N2545,N2549,N2552,
     N2555,N2558,N2561,N2564,N2567,N2570,N2573,N2576,N2579,N2582,
     N2586,N2587,N2588,N2591,N2595,N2599,N2603,N2607,N2611,N2615,
     N2619,N2623,N2627,N2631,N2635,N2639,N2640,N2641,N2644,N2648,
     N2649,N2650,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,
     N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,
     N2671,N2672,N2673,N2674,N2675,N2678,N2682,N2683,N2684,N2687,
     N2690,N2694,N2697,N2700,N2703,N2706,N2709,N2712,N2715,N2718,
     N2721,N2724,N2727,N2731,N2732,N2733,N2736,N2739,N2743,N2744,
     N2745,N2749,N2753,N2757,N2761,N2765,N2769,N2773,N2777,N2781,
     N2785,N2789,N2790,N2791,N2794,N2797,N2801,N2802,N2803,N2806,
     N2807,N2808,N2811,N2812,N2813,N2816,N2817,N2818,N2821,N2822,
     N2823,N2826,N2827,N2828,N2831,N2832,N2833,N2836,N2837,N2838,
     N2841,N2842,N2843,N2846,N2847,N2848,N2851,N2852,N2853,N2856,
     N2857,N2858,N2861,N2864,N2868,N2869,N2870,N2873,N2878,N2881,
     N2884,N2887,N2890,N2893,N2896,N2899,N2902,N2905,N2908,N2912,
     N2913,N2914,N2917,N2921,N2922,N2923,N2926,N2930,N2934,N2938,
     N2942,N2946,N2950,N2954,N2958,N2962,N2966,N2967,N2968,N2971,
     N2975,N2976,N2977,N2980,N2983,N2987,N2988,N2989,N2990,N2991,
     N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
     N3002,N3003,N3004,N3005,N3006,N3007,N3010,N3014,N3015,N3016,
     N3019,N3022,N3026,N3027,N3028,N3031,N3034,N3037,N3040,N3043,
     N3046,N3049,N3052,N3055,N3058,N3062,N3063,N3064,N3067,N3070,
     N3074,N3075,N3076,N3079,N3083,N3087,N3091,N3095,N3099,N3103,
     N3107,N3111,N3115,N3119,N3120,N3121,N3124,N3127,N3131,N3132,
     N3133,N3136,N3140,N3141,N3142,N3145,N3146,N3147,N3150,N3151,
     N3152,N3155,N3156,N3157,N3160,N3161,N3162,N3165,N3166,N3167,
     N3170,N3171,N3172,N3175,N3176,N3177,N3180,N3181,N3182,N3185,
     N3186,N3187,N3190,N3193,N3197,N3198,N3199,N3202,N3206,N3207,
     N3208,N3212,N3215,N3218,N3221,N3224,N3227,N3230,N3233,N3236,
     N3239,N3243,N3244,N3245,N3248,N3252,N3253,N3254,N3257,N3260,
     N3264,N3268,N3272,N3276,N3280,N3284,N3288,N3292,N3296,N3300,
     N3301,N3302,N3305,N3309,N3310,N3311,N3314,N3317,N3321,N3322,
     N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,
     N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3344,
     N3348,N3349,N3350,N3353,N3356,N3360,N3361,N3362,N3365,N3368,
     N3371,N3374,N3377,N3380,N3383,N3386,N3389,N3392,N3396,N3397,
     N3398,N3401,N3404,N3408,N3409,N3410,N3413,N3417,N3421,N3425,
     N3429,N3433,N3437,N3441,N3445,N3449,N3453,N3454,N3455,N3458,
     N3461,N3465,N3466,N3467,N3470,N3474,N3475,N3476,N3479,N3480,
     N3481,N3484,N3485,N3486,N3489,N3490,N3491,N3494,N3495,N3496,
     N3499,N3500,N3501,N3504,N3505,N3506,N3509,N3510,N3511,N3514,
     N3515,N3516,N3519,N3520,N3521,N3524,N3527,N3531,N3532,N3533,
     N3536,N3540,N3541,N3542,N3545,N3548,N3553,N3556,N3559,N3562,
     N3565,N3568,N3571,N3574,N3577,N3581,N3582,N3583,N3586,N3590,
     N3591,N3592,N3595,N3598,N3602,N3603,N3604,N3608,N3612,N3616,
     N3620,N3624,N3628,N3632,N3636,N3637,N3638,N3641,N3645,N3646,
     N3647,N3650,N3653,N3657,N3658,N3659,N3662,N3663,N3664,N3665,
     N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,
     N3676,N3677,N3678,N3681,N3685,N3686,N3687,N3690,N3693,N3697,
     N3698,N3699,N3702,N3706,N3709,N3712,N3715,N3718,N3721,N3724,
     N3727,N3730,N3734,N3735,N3736,N3739,N3742,N3746,N3747,N3748,
     N3751,N3755,N3756,N3757,N3760,N3764,N3768,N3772,N3776,N3780,
     N3784,N3788,N3792,N3793,N3794,N3797,N3800,N3804,N3805,N3806,
     N3809,N3813,N3814,N3815,N3818,N3821,N3825,N3826,N3827,N3830,
     N3831,N3832,N3835,N3836,N3837,N3840,N3841,N3842,N3845,N3846,
     N3847,N3850,N3851,N3852,N3855,N3856,N3857,N3860,N3861,N3862,
     N3865,N3868,N3872,N3873,N3874,N3877,N3881,N3882,N3883,N3886,
     N3889,N3893,N3894,N3896,N3899,N3902,N3905,N3908,N3911,N3914,
     N3917,N3921,N3922,N3923,N3926,N3930,N3931,N3932,N3935,N3938,
     N3942,N3943,N3944,N3947,N3951,N3955,N3959,N3963,N3967,N3971,
     N3975,N3976,N3977,N3980,N3984,N3985,N3986,N3989,N3992,N3996,
     N3997,N3998,N4001,N4005,N4006,N4007,N4008,N4009,N4010,N4011,
     N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4022,N4026,
     N4027,N4028,N4031,N4034,N4038,N4039,N4040,N4043,N4047,N4048,
     N4049,N4052,N4055,N4058,N4061,N4064,N4067,N4070,N4073,N4077,
     N4078,N4079,N4082,N4085,N4089,N4090,N4091,N4094,N4098,N4099,
     N4100,N4103,N4106,N4110,N4114,N4118,N4122,N4126,N4130,N4134,
     N4138,N4139,N4140,N4143,N4146,N4150,N4151,N4152,N4155,N4159,
     N4160,N4161,N4164,N4167,N4171,N4172,N4173,N4174,N4175,N4178,
     N4179,N4180,N4183,N4184,N4185,N4188,N4189,N4190,N4193,N4194,
     N4195,N4198,N4199,N4200,N4203,N4204,N4205,N4208,N4211,N4215,
     N4216,N4217,N4220,N4224,N4225,N4226,N4229,N4232,N4236,N4237,
     N4238,N4242,N4245,N4248,N4251,N4254,N4257,N4260,N4264,N4265,
     N4266,N4269,N4273,N4274,N4275,N4278,N4281,N4285,N4286,N4287,
     N4290,N4294,N4298,N4302,N4306,N4310,N4314,N4318,N4319,N4320,
     N4323,N4327,N4328,N4329,N4332,N4335,N4339,N4340,N4341,N4344,
     N4348,N4349,N4350,N4353,N4354,N4355,N4356,N4357,N4358,N4359,
     N4360,N4361,N4362,N4363,N4364,N4365,N4368,N4372,N4373,N4374,
     N4377,N4380,N4384,N4385,N4386,N4389,N4393,N4394,N4395,N4398,
     N4401,N4405,N4408,N4411,N4414,N4417,N4420,N4423,N4427,N4428,
     N4429,N4432,N4435,N4439,N4440,N4441,N4444,N4448,N4449,N4450,
     N4453,N4456,N4460,N4461,N4462,N4466,N4470,N4474,N4478,N4482,
     N4486,N4487,N4488,N4491,N4494,N4498,N4499,N4500,N4503,N4507,
     N4508,N4509,N4512,N4515,N4519,N4520,N4521,N4524,N4525,N4526,
     N4529,N4530,N4531,N4534,N4535,N4536,N4539,N4540,N4541,N4544,
     N4545,N4546,N4549,N4550,N4551,N4554,N4557,N4561,N4562,N4563,
     N4566,N4570,N4571,N4572,N4575,N4578,N4582,N4583,N4584,N4587,
     N4592,N4595,N4598,N4601,N4604,N4607,N4611,N4612,N4613,N4616,
     N4620,N4621,N4622,N4625,N4628,N4632,N4633,N4634,N4637,N4641,
     N4642,N4643,N4646,N4650,N4654,N4658,N4662,N4666,N4667,N4668,
     N4671,N4675,N4676,N4677,N4680,N4683,N4687,N4688,N4689,N4692,
     N4696,N4697,N4698,N4701,N4704,N4708,N4709,N4710,N4711,N4712,
     N4713,N4714,N4715,N4716,N4717,N4718,N4721,N4725,N4726,N4727,
     N4730,N4733,N4737,N4738,N4739,N4742,N4746,N4747,N4748,N4751,
     N4754,N4758,N4759,N4760,N4763,N4766,N4769,N4772,N4775,N4779,
     N4780,N4781,N4784,N4787,N4791,N4792,N4793,N4796,N4800,N4801,
     N4802,N4805,N4808,N4812,N4813,N4814,N4817,N4821,N4825,N4829,
     N4833,N4837,N4838,N4839,N4842,N4845,N4849,N4850,N4851,N4854,
     N4858,N4859,N4860,N4863,N4866,N4870,N4871,N4872,N4875,N4879,
     N4880,N4881,N4884,N4885,N4886,N4889,N4890,N4891,N4894,N4895,
     N4896,N4899,N4900,N4901,N4904,N4907,N4911,N4912,N4913,N4916,
     N4920,N4921,N4922,N4925,N4928,N4932,N4933,N4934,N4937,N4941,
     N4942,N4943,N4947,N4950,N4953,N4956,N4959,N4963,N4964,N4965,
     N4968,N4972,N4973,N4974,N4977,N4980,N4984,N4985,N4986,N4989,
     N4993,N4994,N4995,N4998,N5001,N5005,N5009,N5013,N5017,N5021,
     N5022,N5023,N5026,N5030,N5031,N5032,N5035,N5038,N5042,N5043,
     N5044,N5047,N5051,N5052,N5053,N5056,N5059,N5063,N5064,N5065,
     N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5076,N5080,
     N5081,N5082,N5085,N5088,N5092,N5093,N5094,N5097,N5101,N5102,
     N5103,N5106,N5109,N5113,N5114,N5115,N5118,N5121,N5124,N5127,
     N5130,N5134,N5135,N5136,N5139,N5142,N5146,N5147,N5148,N5151,
     N5155,N5156,N5157,N5160,N5163,N5167,N5168,N5169,N5172,N5176,
     N5180,N5184,N5188,N5192,N5193,N5194,N5197,N5200,N5204,N5205,
     N5206,N5209,N5213,N5214,N5215,N5218,N5221,N5225,N5226,N5227,
     N5230,N5234,N5235,N5236,N5239,N5240,N5241,N5244,N5245,N5246,
     N5249,N5250,N5251,N5254,N5255,N5256,N5259,N5262,N5266,N5267,
     N5268,N5271,N5275,N5276,N5277,N5280,N5283,N5287,N5288,N5289,
     N5292,N5296,N5297,N5298,N5301,N5304,N5309,N5312,N5315,N5318,
     N5322,N5323,N5324,N5327,N5331,N5332,N5333,N5336,N5339,N5343,
     N5344,N5345,N5348,N5352,N5353,N5354,N5357,N5360,N5364,N5365,
     N5366,N5370,N5374,N5378,N5379,N5380,N5383,N5387,N5388,N5389,
     N5392,N5395,N5399,N5400,N5401,N5404,N5408,N5409,N5410,N5413,
     N5416,N5420,N5421,N5422,N5425,N5426,N5427,N5428,N5429,N5430,
     N5431,N5434,N5438,N5439,N5440,N5443,N5446,N5450,N5451,N5452,
     N5455,N5459,N5460,N5461,N5464,N5467,N5471,N5472,N5473,N5476,
     N5480,N5483,N5486,N5489,N5493,N5494,N5495,N5498,N5501,N5505,
     N5506,N5507,N5510,N5514,N5515,N5516,N5519,N5522,N5526,N5527,
     N5528,N5531,N5535,N5536,N5537,N5540,N5544,N5548,N5552,N5553,
     N5554,N5557,N5560,N5564,N5565,N5566,N5569,N5573,N5574,N5575,
     N5578,N5581,N5585,N5586,N5587,N5590,N5594,N5595,N5596,N5599,
     N5602,N5606,N5607,N5608,N5611,N5612,N5613,N5616,N5617,N5618,
     N5621,N5624,N5628,N5629,N5630,N5633,N5637,N5638,N5639,N5642,
     N5645,N5649,N5650,N5651,N5654,N5658,N5659,N5660,N5663,N5666,
     N5670,N5671,N5673,N5676,N5679,N5683,N5684,N5685,N5688,N5692,
     N5693,N5694,N5697,N5700,N5704,N5705,N5706,N5709,N5713,N5714,
     N5715,N5718,N5721,N5725,N5726,N5727,N5730,N5734,N5738,N5739,
     N5740,N5743,N5747,N5748,N5749,N5752,N5755,N5759,N5760,N5761,
     N5764,N5768,N5769,N5770,N5773,N5776,N5780,N5781,N5782,N5785,
     N5786,N5787,N5788,N5789,N5792,N5796,N5797,N5798,N5801,N5804,
     N5808,N5809,N5810,N5813,N5817,N5818,N5819,N5822,N5825,N5829,
     N5830,N5831,N5834,N5837,N5840,N5844,N5845,N5846,N5849,N5852,
     N5856,N5857,N5858,N5861,N5865,N5866,N5867,N5870,N5873,N5877,
     N5878,N5879,N5882,N5886,N5890,N5891,N5892,N5895,N5898,N5902,
     N5903,N5904,N5907,N5911,N5912,N5913,N5916,N5919,N5923,N5924,
     N5925,N5928,N5929,N5930,N5933,N5934,N5935,N5938,N5941,N5945,
     N5946,N5947,N5950,N5954,N5955,N5956,N5959,N5962,N5966,N5967,
     N5968,N5972,N5975,N5979,N5980,N5981,N5984,N5988,N5989,N5990,
     N5993,N5996,N6000,N6001,N6002,N6005,N6009,N6010,N6011,N6014,
     N6018,N6019,N6020,N6023,N6026,N6030,N6031,N6032,N6035,N6036,
     N6037,N6040,N6044,N6045,N6046,N6049,N6052,N6056,N6057,N6058,
     N6061,N6064,N6068,N6069,N6070,N6073,N6076,N6080,N6081,N6082,
     N6085,N6089,N6090,N6091,N6094,N6097,N6101,N6102,N6103,N6106,
     N6107,N6108,N6111,N6114,N6118,N6119,N6120,N6124,N6128,N6129,
     N6130,N6133,N6134,N6135,N6138,N6141,N6145,N6146,N6147,N6151,
     N6155,N6156,N6157,N6161,N6165,N6166,N6167,N6171,N6175,N6176,
     N6177,N6181,N6185,N6186,N6187,N6191,N6195,N6196,N6197,N6201,
     N6205,N6206,N6207,N6211,N6215,N6216,N6217,N6221,N6225,N6226,
     N6227,N6231,N6235,N6236,N6237,N6241,N6245,N6246,N6247,N6251,
     N6255,N6256,N6257,N6261,N6265,N6266,N6267,N6271,N6275,N6276,
     N6277,N6281,N6285,N6286;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N1_t0,N1_t1,N1_t2,N1_t3,N1_t4,N1_t5,N1_t6,N1_t7,N1_t8,
     N1_t9,N1_t10,N1_t11,N1_t12,N1_t13,N1_t14,N1_t15,N273_t0,N273_t1,N273_t2,
     N273_t3,N273_t4,N273_t5,N273_t6,N273_t7,N273_t8,N273_t9,N273_t10,N273_t11,N273_t12,
     N273_t13,N273_t14,N273_t15,N290_t0,N290_t1,N290_t2,N290_t3,N290_t4,N290_t5,N290_t6,
     N290_t7,N290_t8,N290_t9,N290_t10,N290_t11,N290_t12,N290_t13,N290_t14,N290_t15,N307_t0,
     N307_t1,N307_t2,N307_t3,N307_t4,N307_t5,N307_t6,N307_t7,N307_t8,N307_t9,N307_t10,
     N307_t11,N307_t12,N307_t13,N307_t14,N307_t15,N324_t0,N324_t1,N324_t2,N324_t3,N324_t4,
     N324_t5,N324_t6,N324_t7,N324_t8,N324_t9,N324_t10,N324_t11,N324_t12,N324_t13,N324_t14,
     N324_t15,N341_t0,N341_t1,N341_t2,N341_t3,N341_t4,N341_t5,N341_t6,N341_t7,N341_t8,
     N341_t9,N341_t10,N341_t11,N341_t12,N341_t13,N341_t14,N341_t15,N358_t0,N358_t1,N358_t2,
     N358_t3,N358_t4,N358_t5,N358_t6,N358_t7,N358_t8,N358_t9,N358_t10,N358_t11,N358_t12,
     N358_t13,N358_t14,N358_t15,N375_t0,N375_t1,N375_t2,N375_t3,N375_t4,N375_t5,N375_t6,
     N375_t7,N375_t8,N375_t9,N375_t10,N375_t11,N375_t12,N375_t13,N375_t14,N375_t15,N392_t0,
     N392_t1,N392_t2,N392_t3,N392_t4,N392_t5,N392_t6,N392_t7,N392_t8,N392_t9,N392_t10,
     N392_t11,N392_t12,N392_t13,N392_t14,N392_t15,N409_t0,N409_t1,N409_t2,N409_t3,N409_t4,
     N409_t5,N409_t6,N409_t7,N409_t8,N409_t9,N409_t10,N409_t11,N409_t12,N409_t13,N409_t14,
     N409_t15,N426_t0,N426_t1,N426_t2,N426_t3,N426_t4,N426_t5,N426_t6,N426_t7,N426_t8,
     N426_t9,N426_t10,N426_t11,N426_t12,N426_t13,N426_t14,N426_t15,N443_t0,N443_t1,N443_t2,
     N443_t3,N443_t4,N443_t5,N443_t6,N443_t7,N443_t8,N443_t9,N443_t10,N443_t11,N443_t12,
     N443_t13,N443_t14,N443_t15,N460_t0,N460_t1,N460_t2,N460_t3,N460_t4,N460_t5,N460_t6,
     N460_t7,N460_t8,N460_t9,N460_t10,N460_t11,N460_t12,N460_t13,N460_t14,N460_t15,N477_t0,
     N477_t1,N477_t2,N477_t3,N477_t4,N477_t5,N477_t6,N477_t7,N477_t8,N477_t9,N477_t10,
     N477_t11,N477_t12,N477_t13,N477_t14,N477_t15,N494_t0,N494_t1,N494_t2,N494_t3,N494_t4,
     N494_t5,N494_t6,N494_t7,N494_t8,N494_t9,N494_t10,N494_t11,N494_t12,N494_t13,N494_t14,
     N494_t15,N511_t0,N511_t1,N511_t2,N511_t3,N511_t4,N511_t5,N511_t6,N511_t7,N511_t8,
     N511_t9,N511_t10,N511_t11,N511_t12,N511_t13,N511_t14,N511_t15,N528_t0,N528_t1,N528_t2,
     N528_t3,N528_t4,N528_t5,N528_t6,N528_t7,N528_t8,N528_t9,N528_t10,N528_t11,N528_t12,
     N528_t13,N528_t14,N528_t15,N18_t0,N18_t1,N18_t2,N18_t3,N18_t4,N18_t5,N18_t6,
     N18_t7,N18_t8,N18_t9,N18_t10,N18_t11,N18_t12,N18_t13,N18_t14,N18_t15,N35_t0,
     N35_t1,N35_t2,N35_t3,N35_t4,N35_t5,N35_t6,N35_t7,N35_t8,N35_t9,N35_t10,
     N35_t11,N35_t12,N35_t13,N35_t14,N35_t15,N52_t0,N52_t1,N52_t2,N52_t3,N52_t4,
     N52_t5,N52_t6,N52_t7,N52_t8,N52_t9,N52_t10,N52_t11,N52_t12,N52_t13,N52_t14,
     N52_t15,N69_t0,N69_t1,N69_t2,N69_t3,N69_t4,N69_t5,N69_t6,N69_t7,N69_t8,
     N69_t9,N69_t10,N69_t11,N69_t12,N69_t13,N69_t14,N69_t15,N86_t0,N86_t1,N86_t2,
     N86_t3,N86_t4,N86_t5,N86_t6,N86_t7,N86_t8,N86_t9,N86_t10,N86_t11,N86_t12,
     N86_t13,N86_t14,N86_t15,N103_t0,N103_t1,N103_t2,N103_t3,N103_t4,N103_t5,N103_t6,
     N103_t7,N103_t8,N103_t9,N103_t10,N103_t11,N103_t12,N103_t13,N103_t14,N103_t15,N120_t0,
     N120_t1,N120_t2,N120_t3,N120_t4,N120_t5,N120_t6,N120_t7,N120_t8,N120_t9,N120_t10,
     N120_t11,N120_t12,N120_t13,N120_t14,N120_t15,N137_t0,N137_t1,N137_t2,N137_t3,N137_t4,
     N137_t5,N137_t6,N137_t7,N137_t8,N137_t9,N137_t10,N137_t11,N137_t12,N137_t13,N137_t14,
     N137_t15,N154_t0,N154_t1,N154_t2,N154_t3,N154_t4,N154_t5,N154_t6,N154_t7,N154_t8,
     N154_t9,N154_t10,N154_t11,N154_t12,N154_t13,N154_t14,N154_t15,N171_t0,N171_t1,N171_t2,
     N171_t3,N171_t4,N171_t5,N171_t6,N171_t7,N171_t8,N171_t9,N171_t10,N171_t11,N171_t12,
     N171_t13,N171_t14,N171_t15,N188_t0,N188_t1,N188_t2,N188_t3,N188_t4,N188_t5,N188_t6,
     N188_t7,N188_t8,N188_t9,N188_t10,N188_t11,N188_t12,N188_t13,N188_t14,N188_t15,N205_t0,
     N205_t1,N205_t2,N205_t3,N205_t4,N205_t5,N205_t6,N205_t7,N205_t8,N205_t9,N205_t10,
     N205_t11,N205_t12,N205_t13,N205_t14,N205_t15,N222_t0,N222_t1,N222_t2,N222_t3,N222_t4,
     N222_t5,N222_t6,N222_t7,N222_t8,N222_t9,N222_t10,N222_t11,N222_t12,N222_t13,N222_t14,
     N222_t15,N239_t0,N239_t1,N239_t2,N239_t3,N239_t4,N239_t5,N239_t6,N239_t7,N239_t8,
     N239_t9,N239_t10,N239_t11,N239_t12,N239_t13,N239_t14,N239_t15,N256_t0,N256_t1,N256_t2,
     N256_t3,N256_t4,N256_t5,N256_t6,N256_t7,N256_t8,N256_t9,N256_t10,N256_t11,N256_t12,
     N256_t13,N256_t14,N256_t15,N591_t0,N591_t1,N639_t0,N639_t1,N687_t0,N687_t1,N735_t0,
     N735_t1,N783_t0,N783_t1,N831_t0,N831_t1,N879_t0,N879_t1,N927_t0,N927_t1,N975_t0,
     N975_t1,N1023_t0,N1023_t1,N1071_t0,N1071_t1,N1119_t0,N1119_t1,N1167_t0,N1167_t1,N1215_t0,
     N1215_t1,N1263_t0,N1263_t1,N1311_t0,N1311_t1,N1311_t2,N1315_t0,N1315_t1,N1315_t2,N1319_t0,
     N1319_t1,N1319_t2,N1323_t0,N1323_t1,N1323_t2,N1327_t0,N1327_t1,N1327_t2,N1331_t0,N1331_t1,
     N1331_t2,N1335_t0,N1335_t1,N1335_t2,N1339_t0,N1339_t1,N1339_t2,N1343_t0,N1343_t1,N1343_t2,
     N1347_t0,N1347_t1,N1347_t2,N1351_t0,N1351_t1,N1351_t2,N1355_t0,N1355_t1,N1355_t2,N1359_t0,
     N1359_t1,N1359_t2,N1363_t0,N1363_t1,N1363_t2,N1367_t0,N1367_t1,N1367_t2,N1401_t0,N1401_t1,
     N546_t0,N546_t1,N1404_t0,N1404_t1,N594_t0,N594_t1,N1407_t0,N1407_t1,N642_t0,N642_t1,
     N1410_t0,N1410_t1,N690_t0,N690_t1,N1413_t0,N1413_t1,N738_t0,N738_t1,N1416_t0,N1416_t1,
     N786_t0,N786_t1,N1419_t0,N1419_t1,N834_t0,N834_t1,N1422_t0,N1422_t1,N882_t0,N882_t1,
     N1425_t0,N1425_t1,N930_t0,N930_t1,N1428_t0,N1428_t1,N978_t0,N978_t1,N1431_t0,N1431_t1,
     N1026_t0,N1026_t1,N1434_t0,N1434_t1,N1074_t0,N1074_t1,N1437_t0,N1437_t1,N1122_t0,N1122_t1,
     N1440_t0,N1440_t1,N1170_t0,N1170_t1,N1443_t0,N1443_t1,N1218_t0,N1218_t1,N1446_t0,N1446_t1,
     N1446_t2,N1450_t0,N1450_t1,N1450_t2,N1454_t0,N1454_t1,N1454_t2,N1458_t0,N1458_t1,N1458_t2,
     N1462_t0,N1462_t1,N1462_t2,N1466_t0,N1466_t1,N1466_t2,N1470_t0,N1470_t1,N1470_t2,N1474_t0,
     N1474_t1,N1474_t2,N1478_t0,N1478_t1,N1478_t2,N1482_t0,N1482_t1,N1482_t2,N1486_t0,N1486_t1,
     N1486_t2,N1490_t0,N1490_t1,N1490_t2,N1494_t0,N1494_t1,N1494_t2,N1498_t0,N1498_t1,N1498_t2,
     N1502_t0,N1502_t1,N1502_t2,N1266_t0,N1266_t1,N1578_t0,N1578_t1,N1582_t0,N1582_t1,N1508_t0,
     N1508_t1,N1585_t0,N1585_t1,N1513_t0,N1513_t1,N1588_t0,N1588_t1,N1518_t0,N1518_t1,N1591_t0,
     N1591_t1,N1523_t0,N1523_t1,N1594_t0,N1594_t1,N1528_t0,N1528_t1,N1597_t0,N1597_t1,N1533_t0,
     N1533_t1,N1600_t0,N1600_t1,N1538_t0,N1538_t1,N1603_t0,N1603_t1,N1543_t0,N1543_t1,N1606_t0,
     N1606_t1,N1548_t0,N1548_t1,N1609_t0,N1609_t1,N1553_t0,N1553_t1,N1612_t0,N1612_t1,N1558_t0,
     N1558_t1,N1615_t0,N1615_t1,N1563_t0,N1563_t1,N1618_t0,N1618_t1,N1568_t0,N1568_t1,N1621_t0,
     N1621_t1,N1573_t0,N1573_t1,N1624_t0,N1624_t1,N1624_t2,N1628_t0,N1628_t1,N1628_t2,N1632_t0,
     N1632_t1,N1632_t2,N1636_t0,N1636_t1,N1636_t2,N1640_t0,N1640_t1,N1640_t2,N1644_t0,N1644_t1,
     N1644_t2,N1648_t0,N1648_t1,N1648_t2,N1652_t0,N1652_t1,N1652_t2,N1656_t0,N1656_t1,N1656_t2,
     N1660_t0,N1660_t1,N1660_t2,N1664_t0,N1664_t1,N1664_t2,N1668_t0,N1668_t1,N1668_t2,N1672_t0,
     N1672_t1,N1672_t2,N1676_t0,N1676_t1,N1676_t2,N1680_t0,N1680_t1,N1680_t2,N1714_t0,N1714_t1,
     N1221_t0,N1221_t1,N1717_t0,N1717_t1,N549_t0,N549_t1,N1720_t0,N1720_t1,N597_t0,N597_t1,
     N1723_t0,N1723_t1,N645_t0,N645_t1,N1726_t0,N1726_t1,N693_t0,N693_t1,N1729_t0,N1729_t1,
     N741_t0,N741_t1,N1732_t0,N1732_t1,N789_t0,N789_t1,N1735_t0,N1735_t1,N837_t0,N837_t1,
     N1738_t0,N1738_t1,N885_t0,N885_t1,N1741_t0,N1741_t1,N933_t0,N933_t1,N1744_t0,N1744_t1,
     N981_t0,N981_t1,N1747_t0,N1747_t1,N1029_t0,N1029_t1,N1750_t0,N1750_t1,N1077_t0,N1077_t1,
     N1753_t0,N1753_t1,N1125_t0,N1125_t1,N1756_t0,N1756_t1,N1173_t0,N1173_t1,N1759_t0,N1759_t1,
     N1759_t2,N1763_t0,N1763_t1,N1763_t2,N1767_t0,N1767_t1,N1767_t2,N1771_t0,N1771_t1,N1771_t2,
     N1775_t0,N1775_t1,N1775_t2,N1779_t0,N1779_t1,N1779_t2,N1783_t0,N1783_t1,N1783_t2,N1787_t0,
     N1787_t1,N1787_t2,N1791_t0,N1791_t1,N1791_t2,N1795_t0,N1795_t1,N1795_t2,N1799_t0,N1799_t1,
     N1799_t2,N1803_t0,N1803_t1,N1803_t2,N1807_t0,N1807_t1,N1807_t2,N1811_t0,N1811_t1,N1811_t2,
     N1815_t0,N1815_t1,N1815_t2,N1269_t0,N1269_t1,N1821_t0,N1821_t1,N1894_t0,N1894_t1,N1891_t0,
     N1891_t1,N1897_t0,N1897_t1,N1897_t2,N1902_t0,N1902_t1,N1826_t0,N1826_t1,N1905_t0,N1905_t1,
     N1831_t0,N1831_t1,N1908_t0,N1908_t1,N1836_t0,N1836_t1,N1911_t0,N1911_t1,N1841_t0,N1841_t1,
     N1914_t0,N1914_t1,N1846_t0,N1846_t1,N1917_t0,N1917_t1,N1851_t0,N1851_t1,N1920_t0,N1920_t1,
     N1856_t0,N1856_t1,N1923_t0,N1923_t1,N1861_t0,N1861_t1,N1926_t0,N1926_t1,N1866_t0,N1866_t1,
     N1929_t0,N1929_t1,N1871_t0,N1871_t1,N1932_t0,N1932_t1,N1876_t0,N1876_t1,N1935_t0,N1935_t1,
     N1881_t0,N1881_t1,N1938_t0,N1938_t1,N1886_t0,N1886_t1,N1941_t0,N1941_t1,N1941_t2,N1947_t0,
     N1947_t1,N1947_t2,N1951_t0,N1951_t1,N1951_t2,N1955_t0,N1955_t1,N1955_t2,N1959_t0,N1959_t1,
     N1959_t2,N1963_t0,N1963_t1,N1963_t2,N1967_t0,N1967_t1,N1967_t2,N1971_t0,N1971_t1,N1971_t2,
     N1975_t0,N1975_t1,N1975_t2,N1979_t0,N1979_t1,N1979_t2,N1983_t0,N1983_t1,N1983_t2,N1987_t0,
     N1987_t1,N1987_t2,N1991_t0,N1991_t1,N1991_t2,N1995_t0,N1995_t1,N1995_t2,N2001_t0,N2001_t1,
     N1224_t0,N1224_t1,N2030_t0,N2030_t1,N1176_t0,N1176_t1,N2033_t0,N2033_t1,N2033_t2,N2037_t0,
     N2037_t1,N552_t0,N552_t1,N2040_t0,N2040_t1,N600_t0,N600_t1,N2043_t0,N2043_t1,N648_t0,
     N648_t1,N2046_t0,N2046_t1,N696_t0,N696_t1,N2049_t0,N2049_t1,N744_t0,N744_t1,N2052_t0,
     N2052_t1,N792_t0,N792_t1,N2055_t0,N2055_t1,N840_t0,N840_t1,N2058_t0,N2058_t1,N888_t0,
     N888_t1,N2061_t0,N2061_t1,N936_t0,N936_t1,N2064_t0,N2064_t1,N984_t0,N984_t1,N2067_t0,
     N2067_t1,N1032_t0,N1032_t1,N2070_t0,N2070_t1,N1080_t0,N1080_t1,N2073_t0,N2073_t1,N1128_t0,
     N1128_t1,N2076_t0,N2076_t1,N2076_t2,N1272_t0,N1272_t1,N2082_t0,N2082_t1,N2085_t0,N2085_t1,
     N2085_t2,N2089_t0,N2089_t1,N2089_t2,N2093_t0,N2093_t1,N2093_t2,N2097_t0,N2097_t1,N2097_t2,
     N2101_t0,N2101_t1,N2101_t2,N2105_t0,N2105_t1,N2105_t2,N2109_t0,N2109_t1,N2109_t2,N2113_t0,
     N2113_t1,N2113_t2,N2117_t0,N2117_t1,N2117_t2,N2121_t0,N2121_t1,N2121_t2,N2125_t0,N2125_t1,
     N2125_t2,N2129_t0,N2129_t1,N2129_t2,N2133_t0,N2133_t1,N2133_t2,N2142_t0,N2142_t1,N2139_t0,
     N2139_t1,N2145_t0,N2145_t1,N2145_t2,N2214_t0,N2214_t1,N2211_t0,N2211_t1,N2217_t0,N2217_t1,
     N2217_t2,N2224_t0,N2224_t1,N2151_t0,N2151_t1,N2227_t0,N2227_t1,N2156_t0,N2156_t1,N2230_t0,
     N2230_t1,N2161_t0,N2161_t1,N2233_t0,N2233_t1,N2166_t0,N2166_t1,N2236_t0,N2236_t1,N2171_t0,
     N2171_t1,N2239_t0,N2239_t1,N2176_t0,N2176_t1,N2242_t0,N2242_t1,N2181_t0,N2181_t1,N2245_t0,
     N2245_t1,N2186_t0,N2186_t1,N2248_t0,N2248_t1,N2191_t0,N2191_t1,N2251_t0,N2251_t1,N2196_t0,
     N2196_t1,N2254_t0,N2254_t1,N2201_t0,N2201_t1,N2257_t0,N2257_t1,N2206_t0,N2206_t1,N2260_t0,
     N2260_t1,N2260_t2,N2266_t0,N2266_t1,N1227_t0,N1227_t1,N2269_t0,N2269_t1,N2269_t2,N2273_t0,
     N2273_t1,N2273_t2,N2277_t0,N2277_t1,N2277_t2,N2281_t0,N2281_t1,N2281_t2,N2285_t0,N2285_t1,
     N2285_t2,N2289_t0,N2289_t1,N2289_t2,N2293_t0,N2293_t1,N2293_t2,N2297_t0,N2297_t1,N2297_t2,
     N2301_t0,N2301_t1,N2301_t2,N2305_t0,N2305_t1,N2305_t2,N2309_t0,N2309_t1,N2309_t2,N2313_t0,
     N2313_t1,N2313_t2,N2319_t0,N2319_t1,N1179_t0,N1179_t1,N2322_t0,N2322_t1,N2322_t2,N2350_t0,
     N2350_t1,N1131_t0,N1131_t1,N2353_t0,N2353_t1,N2353_t2,N1275_t0,N1275_t1,N2359_t0,N2359_t1,
     N2362_t0,N2362_t1,N555_t0,N555_t1,N2365_t0,N2365_t1,N603_t0,N603_t1,N2368_t0,N2368_t1,
     N651_t0,N651_t1,N2371_t0,N2371_t1,N699_t0,N699_t1,N2374_t0,N2374_t1,N747_t0,N747_t1,
     N2377_t0,N2377_t1,N795_t0,N795_t1,N2380_t0,N2380_t1,N843_t0,N843_t1,N2383_t0,N2383_t1,
     N891_t0,N891_t1,N2386_t0,N2386_t1,N939_t0,N939_t1,N2389_t0,N2389_t1,N987_t0,N987_t1,
     N2392_t0,N2392_t1,N1035_t0,N1035_t1,N2395_t0,N2395_t1,N1083_t0,N1083_t1,N2398_t0,N2398_t1,
     N2398_t2,N2407_t0,N2407_t1,N2404_t0,N2404_t1,N2410_t0,N2410_t1,N2410_t2,N2414_t0,N2414_t1,
     N2414_t2,N2418_t0,N2418_t1,N2418_t2,N2422_t0,N2422_t1,N2422_t2,N2426_t0,N2426_t1,N2426_t2,
     N2430_t0,N2430_t1,N2430_t2,N2434_t0,N2434_t1,N2434_t2,N2438_t0,N2438_t1,N2438_t2,N2442_t0,
     N2442_t1,N2442_t2,N2446_t0,N2446_t1,N2446_t2,N2450_t0,N2450_t1,N2450_t2,N2454_t0,N2454_t1,
     N2454_t2,N2458_t0,N2458_t1,N2458_t2,N2467_t0,N2467_t1,N2464_t0,N2464_t1,N2470_t0,N2470_t1,
     N2470_t2,N2536_t0,N2536_t1,N2533_t0,N2533_t1,N2539_t0,N2539_t1,N2539_t2,N2545_t0,N2545_t1,
     N1230_t0,N1230_t1,N2549_t0,N2549_t1,N2478_t0,N2478_t1,N2552_t0,N2552_t1,N2483_t0,N2483_t1,
     N2555_t0,N2555_t1,N2488_t0,N2488_t1,N2558_t0,N2558_t1,N2493_t0,N2493_t1,N2561_t0,N2561_t1,
     N2498_t0,N2498_t1,N2564_t0,N2564_t1,N2503_t0,N2503_t1,N2567_t0,N2567_t1,N2508_t0,N2508_t1,
     N2570_t0,N2570_t1,N2513_t0,N2513_t1,N2573_t0,N2573_t1,N2518_t0,N2518_t1,N2576_t0,N2576_t1,
     N2523_t0,N2523_t1,N2579_t0,N2579_t1,N2528_t0,N2528_t1,N2582_t0,N2582_t1,N2582_t2,N2588_t0,
     N2588_t1,N1182_t0,N1182_t1,N2591_t0,N2591_t1,N2591_t2,N2595_t0,N2595_t1,N2595_t2,N2599_t0,
     N2599_t1,N2599_t2,N2603_t0,N2603_t1,N2603_t2,N2607_t0,N2607_t1,N2607_t2,N2611_t0,N2611_t1,
     N2611_t2,N2615_t0,N2615_t1,N2615_t2,N2619_t0,N2619_t1,N2619_t2,N2623_t0,N2623_t1,N2623_t2,
     N2627_t0,N2627_t1,N2627_t2,N2631_t0,N2631_t1,N2631_t2,N2635_t0,N2635_t1,N2635_t2,N2641_t0,
     N2641_t1,N1134_t0,N1134_t1,N2644_t0,N2644_t1,N2644_t2,N1278_t0,N1278_t1,N2650_t0,N2650_t1,
     N2675_t0,N2675_t1,N1086_t0,N1086_t1,N2678_t0,N2678_t1,N2678_t2,N2687_t0,N2687_t1,N2684_t0,
     N2684_t1,N2690_t0,N2690_t1,N2690_t2,N2694_t0,N2694_t1,N558_t0,N558_t1,N2697_t0,N2697_t1,
     N606_t0,N606_t1,N2700_t0,N2700_t1,N654_t0,N654_t1,N2703_t0,N2703_t1,N702_t0,N702_t1,
     N2706_t0,N2706_t1,N750_t0,N750_t1,N2709_t0,N2709_t1,N798_t0,N798_t1,N2712_t0,N2712_t1,
     N846_t0,N846_t1,N2715_t0,N2715_t1,N894_t0,N894_t1,N2718_t0,N2718_t1,N942_t0,N942_t1,
     N2721_t0,N2721_t1,N990_t0,N990_t1,N2724_t0,N2724_t1,N1038_t0,N1038_t1,N2727_t0,N2727_t1,
     N2727_t2,N2736_t0,N2736_t1,N2733_t0,N2733_t1,N2739_t0,N2739_t1,N2739_t2,N2745_t0,N2745_t1,
     N2745_t2,N2749_t0,N2749_t1,N2749_t2,N2753_t0,N2753_t1,N2753_t2,N2757_t0,N2757_t1,N2757_t2,
     N2761_t0,N2761_t1,N2761_t2,N2765_t0,N2765_t1,N2765_t2,N2769_t0,N2769_t1,N2769_t2,N2773_t0,
     N2773_t1,N2773_t2,N2777_t0,N2777_t1,N2777_t2,N2781_t0,N2781_t1,N2781_t2,N2785_t0,N2785_t1,
     N2785_t2,N2794_t0,N2794_t1,N2791_t0,N2791_t1,N2797_t0,N2797_t1,N2797_t2,N2803_t0,N2803_t1,
     N1233_t0,N1233_t1,N2861_t0,N2861_t1,N2858_t0,N2858_t1,N2864_t0,N2864_t1,N2864_t2,N2870_t0,
     N2870_t1,N1185_t0,N1185_t1,N2873_t0,N2873_t1,N2873_t2,N2878_t0,N2878_t1,N2808_t0,N2808_t1,
     N2881_t0,N2881_t1,N2813_t0,N2813_t1,N2884_t0,N2884_t1,N2818_t0,N2818_t1,N2887_t0,N2887_t1,
     N2823_t0,N2823_t1,N2890_t0,N2890_t1,N2828_t0,N2828_t1,N2893_t0,N2893_t1,N2833_t0,N2833_t1,
     N2896_t0,N2896_t1,N2838_t0,N2838_t1,N2899_t0,N2899_t1,N2843_t0,N2843_t1,N2902_t0,N2902_t1,
     N2848_t0,N2848_t1,N2905_t0,N2905_t1,N2853_t0,N2853_t1,N2908_t0,N2908_t1,N2908_t2,N2914_t0,
     N2914_t1,N1137_t0,N1137_t1,N2917_t0,N2917_t1,N2917_t2,N1281_t0,N1281_t1,N2923_t0,N2923_t1,
     N2926_t0,N2926_t1,N2926_t2,N2930_t0,N2930_t1,N2930_t2,N2934_t0,N2934_t1,N2934_t2,N2938_t0,
     N2938_t1,N2938_t2,N2942_t0,N2942_t1,N2942_t2,N2946_t0,N2946_t1,N2946_t2,N2950_t0,N2950_t1,
     N2950_t2,N2954_t0,N2954_t1,N2954_t2,N2958_t0,N2958_t1,N2958_t2,N2962_t0,N2962_t1,N2962_t2,
     N2968_t0,N2968_t1,N1089_t0,N1089_t1,N2971_t0,N2971_t1,N2971_t2,N2980_t0,N2980_t1,N2977_t0,
     N2977_t1,N2983_t0,N2983_t1,N2983_t2,N3007_t0,N3007_t1,N1041_t0,N1041_t1,N3010_t0,N3010_t1,
     N3010_t2,N3019_t0,N3019_t1,N3016_t0,N3016_t1,N3022_t0,N3022_t1,N3022_t2,N3028_t0,N3028_t1,
     N561_t0,N561_t1,N3031_t0,N3031_t1,N609_t0,N609_t1,N3034_t0,N3034_t1,N657_t0,N657_t1,
     N3037_t0,N3037_t1,N705_t0,N705_t1,N3040_t0,N3040_t1,N753_t0,N753_t1,N3043_t0,N3043_t1,
     N801_t0,N801_t1,N3046_t0,N3046_t1,N849_t0,N849_t1,N3049_t0,N3049_t1,N897_t0,N897_t1,
     N3052_t0,N3052_t1,N945_t0,N945_t1,N3055_t0,N3055_t1,N993_t0,N993_t1,N3058_t0,N3058_t1,
     N3058_t2,N3067_t0,N3067_t1,N3064_t0,N3064_t1,N3070_t0,N3070_t1,N3070_t2,N3076_t0,N3076_t1,
     N1236_t0,N1236_t1,N3079_t0,N3079_t1,N3079_t2,N3083_t0,N3083_t1,N3083_t2,N3087_t0,N3087_t1,
     N3087_t2,N3091_t0,N3091_t1,N3091_t2,N3095_t0,N3095_t1,N3095_t2,N3099_t0,N3099_t1,N3099_t2,
     N3103_t0,N3103_t1,N3103_t2,N3107_t0,N3107_t1,N3107_t2,N3111_t0,N3111_t1,N3111_t2,N3115_t0,
     N3115_t1,N3115_t2,N3124_t0,N3124_t1,N3121_t0,N3121_t1,N3127_t0,N3127_t1,N3127_t2,N3133_t0,
     N3133_t1,N1188_t0,N1188_t1,N3136_t0,N3136_t1,N3136_t2,N3190_t0,N3190_t1,N3187_t0,N3187_t1,
     N3193_t0,N3193_t1,N3193_t2,N3199_t0,N3199_t1,N1140_t0,N1140_t1,N3202_t0,N3202_t1,N3202_t2,
     N1284_t0,N1284_t1,N3208_t0,N3208_t1,N3212_t0,N3212_t1,N3142_t0,N3142_t1,N3215_t0,N3215_t1,
     N3147_t0,N3147_t1,N3218_t0,N3218_t1,N3152_t0,N3152_t1,N3221_t0,N3221_t1,N3157_t0,N3157_t1,
     N3224_t0,N3224_t1,N3162_t0,N3162_t1,N3227_t0,N3227_t1,N3167_t0,N3167_t1,N3230_t0,N3230_t1,
     N3172_t0,N3172_t1,N3233_t0,N3233_t1,N3177_t0,N3177_t1,N3236_t0,N3236_t1,N3182_t0,N3182_t1,
     N3239_t0,N3239_t1,N3239_t2,N3245_t0,N3245_t1,N1092_t0,N1092_t1,N3248_t0,N3248_t1,N3248_t2,
     N3257_t0,N3257_t1,N3254_t0,N3254_t1,N3260_t0,N3260_t1,N3260_t2,N3264_t0,N3264_t1,N3264_t2,
     N3268_t0,N3268_t1,N3268_t2,N3272_t0,N3272_t1,N3272_t2,N3276_t0,N3276_t1,N3276_t2,N3280_t0,
     N3280_t1,N3280_t2,N3284_t0,N3284_t1,N3284_t2,N3288_t0,N3288_t1,N3288_t2,N3292_t0,N3292_t1,
     N3292_t2,N3296_t0,N3296_t1,N3296_t2,N3302_t0,N3302_t1,N1044_t0,N1044_t1,N3305_t0,N3305_t1,
     N3305_t2,N3314_t0,N3314_t1,N3311_t0,N3311_t1,N3317_t0,N3317_t1,N3317_t2,N3341_t0,N3341_t1,
     N996_t0,N996_t1,N3344_t0,N3344_t1,N3344_t2,N3353_t0,N3353_t1,N3350_t0,N3350_t1,N3356_t0,
     N3356_t1,N3356_t2,N3362_t0,N3362_t1,N1239_t0,N1239_t1,N3365_t0,N3365_t1,N564_t0,N564_t1,
     N3368_t0,N3368_t1,N612_t0,N612_t1,N3371_t0,N3371_t1,N660_t0,N660_t1,N3374_t0,N3374_t1,
     N708_t0,N708_t1,N3377_t0,N3377_t1,N756_t0,N756_t1,N3380_t0,N3380_t1,N804_t0,N804_t1,
     N3383_t0,N3383_t1,N852_t0,N852_t1,N3386_t0,N3386_t1,N900_t0,N900_t1,N3389_t0,N3389_t1,
     N948_t0,N948_t1,N3392_t0,N3392_t1,N3392_t2,N3401_t0,N3401_t1,N3398_t0,N3398_t1,N3404_t0,
     N3404_t1,N3404_t2,N3410_t0,N3410_t1,N1191_t0,N1191_t1,N3413_t0,N3413_t1,N3413_t2,N3417_t0,
     N3417_t1,N3417_t2,N3421_t0,N3421_t1,N3421_t2,N3425_t0,N3425_t1,N3425_t2,N3429_t0,N3429_t1,
     N3429_t2,N3433_t0,N3433_t1,N3433_t2,N3437_t0,N3437_t1,N3437_t2,N3441_t0,N3441_t1,N3441_t2,
     N3445_t0,N3445_t1,N3445_t2,N3449_t0,N3449_t1,N3449_t2,N3458_t0,N3458_t1,N3455_t0,N3455_t1,
     N3461_t0,N3461_t1,N3461_t2,N3467_t0,N3467_t1,N1143_t0,N1143_t1,N3470_t0,N3470_t1,N3470_t2,
     N1287_t0,N1287_t1,N3476_t0,N3476_t1,N3524_t0,N3524_t1,N3521_t0,N3521_t1,N3527_t0,N3527_t1,
     N3527_t2,N3533_t0,N3533_t1,N1095_t0,N1095_t1,N3536_t0,N3536_t1,N3536_t2,N3545_t0,N3545_t1,
     N3542_t0,N3542_t1,N3548_t0,N3548_t1,N3548_t2,N3553_t0,N3553_t1,N3481_t0,N3481_t1,N3556_t0,
     N3556_t1,N3486_t0,N3486_t1,N3559_t0,N3559_t1,N3491_t0,N3491_t1,N3562_t0,N3562_t1,N3496_t0,
     N3496_t1,N3565_t0,N3565_t1,N3501_t0,N3501_t1,N3568_t0,N3568_t1,N3506_t0,N3506_t1,N3571_t0,
     N3571_t1,N3511_t0,N3511_t1,N3574_t0,N3574_t1,N3516_t0,N3516_t1,N3577_t0,N3577_t1,N3577_t2,
     N3583_t0,N3583_t1,N1047_t0,N1047_t1,N3586_t0,N3586_t1,N3586_t2,N3595_t0,N3595_t1,N3592_t0,
     N3592_t1,N3598_t0,N3598_t1,N3598_t2,N3604_t0,N3604_t1,N3604_t2,N3608_t0,N3608_t1,N3608_t2,
     N3612_t0,N3612_t1,N3612_t2,N3616_t0,N3616_t1,N3616_t2,N3620_t0,N3620_t1,N3620_t2,N3624_t0,
     N3624_t1,N3624_t2,N3628_t0,N3628_t1,N3628_t2,N3632_t0,N3632_t1,N3632_t2,N3638_t0,N3638_t1,
     N999_t0,N999_t1,N3641_t0,N3641_t1,N3641_t2,N3650_t0,N3650_t1,N3647_t0,N3647_t1,N3653_t0,
     N3653_t1,N3653_t2,N3659_t0,N3659_t1,N1242_t0,N1242_t1,N3678_t0,N3678_t1,N951_t0,N951_t1,
     N3681_t0,N3681_t1,N3681_t2,N3690_t0,N3690_t1,N3687_t0,N3687_t1,N3693_t0,N3693_t1,N3693_t2,
     N3699_t0,N3699_t1,N1194_t0,N1194_t1,N3702_t0,N3702_t1,N3702_t2,N3706_t0,N3706_t1,N567_t0,
     N567_t1,N3709_t0,N3709_t1,N615_t0,N615_t1,N3712_t0,N3712_t1,N663_t0,N663_t1,N3715_t0,
     N3715_t1,N711_t0,N711_t1,N3718_t0,N3718_t1,N759_t0,N759_t1,N3721_t0,N3721_t1,N807_t0,
     N807_t1,N3724_t0,N3724_t1,N855_t0,N855_t1,N3727_t0,N3727_t1,N903_t0,N903_t1,N3730_t0,
     N3730_t1,N3730_t2,N3739_t0,N3739_t1,N3736_t0,N3736_t1,N3742_t0,N3742_t1,N3742_t2,N3748_t0,
     N3748_t1,N1146_t0,N1146_t1,N3751_t0,N3751_t1,N3751_t2,N1290_t0,N1290_t1,N3757_t0,N3757_t1,
     N3760_t0,N3760_t1,N3760_t2,N3764_t0,N3764_t1,N3764_t2,N3768_t0,N3768_t1,N3768_t2,N3772_t0,
     N3772_t1,N3772_t2,N3776_t0,N3776_t1,N3776_t2,N3780_t0,N3780_t1,N3780_t2,N3784_t0,N3784_t1,
     N3784_t2,N3788_t0,N3788_t1,N3788_t2,N3797_t0,N3797_t1,N3794_t0,N3794_t1,N3800_t0,N3800_t1,
     N3800_t2,N3806_t0,N3806_t1,N1098_t0,N1098_t1,N3809_t0,N3809_t1,N3809_t2,N3818_t0,N3818_t1,
     N3815_t0,N3815_t1,N3821_t0,N3821_t1,N3821_t2,N3865_t0,N3865_t1,N3862_t0,N3862_t1,N3868_t0,
     N3868_t1,N3868_t2,N3874_t0,N3874_t1,N1050_t0,N1050_t1,N3877_t0,N3877_t1,N3877_t2,N3886_t0,
     N3886_t1,N3883_t0,N3883_t1,N3889_t0,N3889_t1,N3889_t2,N3896_t0,N3896_t1,N3827_t0,N3827_t1,
     N3899_t0,N3899_t1,N3832_t0,N3832_t1,N3902_t0,N3902_t1,N3837_t0,N3837_t1,N3905_t0,N3905_t1,
     N3842_t0,N3842_t1,N3908_t0,N3908_t1,N3847_t0,N3847_t1,N3911_t0,N3911_t1,N3852_t0,N3852_t1,
     N3914_t0,N3914_t1,N3857_t0,N3857_t1,N3917_t0,N3917_t1,N3917_t2,N3923_t0,N3923_t1,N1002_t0,
     N1002_t1,N3926_t0,N3926_t1,N3926_t2,N3935_t0,N3935_t1,N3932_t0,N3932_t1,N3938_t0,N3938_t1,
     N3938_t2,N3944_t0,N3944_t1,N1245_t0,N1245_t1,N3947_t0,N3947_t1,N3947_t2,N3951_t0,N3951_t1,
     N3951_t2,N3955_t0,N3955_t1,N3955_t2,N3959_t0,N3959_t1,N3959_t2,N3963_t0,N3963_t1,N3963_t2,
     N3967_t0,N3967_t1,N3967_t2,N3971_t0,N3971_t1,N3971_t2,N3977_t0,N3977_t1,N954_t0,N954_t1,
     N3980_t0,N3980_t1,N3980_t2,N3989_t0,N3989_t1,N3986_t0,N3986_t1,N3992_t0,N3992_t1,N3992_t2,
     N3998_t0,N3998_t1,N1197_t0,N1197_t1,N4001_t0,N4001_t1,N4001_t2,N4019_t0,N4019_t1,N906_t0,
     N906_t1,N4022_t0,N4022_t1,N4022_t2,N4031_t0,N4031_t1,N4028_t0,N4028_t1,N4034_t0,N4034_t1,
     N4034_t2,N4040_t0,N4040_t1,N1149_t0,N1149_t1,N4043_t0,N4043_t1,N4043_t2,N1293_t0,N1293_t1,
     N4049_t0,N4049_t1,N4052_t0,N4052_t1,N570_t0,N570_t1,N4055_t0,N4055_t1,N618_t0,N618_t1,
     N4058_t0,N4058_t1,N666_t0,N666_t1,N4061_t0,N4061_t1,N714_t0,N714_t1,N4064_t0,N4064_t1,
     N762_t0,N762_t1,N4067_t0,N4067_t1,N810_t0,N810_t1,N4070_t0,N4070_t1,N858_t0,N858_t1,
     N4073_t0,N4073_t1,N4073_t2,N4082_t0,N4082_t1,N4079_t0,N4079_t1,N4085_t0,N4085_t1,N4085_t2,
     N4091_t0,N4091_t1,N1101_t0,N1101_t1,N4094_t0,N4094_t1,N4094_t2,N4103_t0,N4103_t1,N4100_t0,
     N4100_t1,N4106_t0,N4106_t1,N4106_t2,N4110_t0,N4110_t1,N4110_t2,N4114_t0,N4114_t1,N4114_t2,
     N4118_t0,N4118_t1,N4118_t2,N4122_t0,N4122_t1,N4122_t2,N4126_t0,N4126_t1,N4126_t2,N4130_t0,
     N4130_t1,N4130_t2,N4134_t0,N4134_t1,N4134_t2,N4143_t0,N4143_t1,N4140_t0,N4140_t1,N4146_t0,
     N4146_t1,N4146_t2,N4152_t0,N4152_t1,N1053_t0,N1053_t1,N4155_t0,N4155_t1,N4155_t2,N4164_t0,
     N4164_t1,N4161_t0,N4161_t1,N4167_t0,N4167_t1,N4167_t2,N4208_t0,N4208_t1,N4205_t0,N4205_t1,
     N4211_t0,N4211_t1,N4211_t2,N4217_t0,N4217_t1,N1005_t0,N1005_t1,N4220_t0,N4220_t1,N4220_t2,
     N4229_t0,N4229_t1,N4226_t0,N4226_t1,N4232_t0,N4232_t1,N4232_t2,N4238_t0,N4238_t1,N1248_t0,
     N1248_t1,N4242_t0,N4242_t1,N4175_t0,N4175_t1,N4245_t0,N4245_t1,N4180_t0,N4180_t1,N4248_t0,
     N4248_t1,N4185_t0,N4185_t1,N4251_t0,N4251_t1,N4190_t0,N4190_t1,N4254_t0,N4254_t1,N4195_t0,
     N4195_t1,N4257_t0,N4257_t1,N4200_t0,N4200_t1,N4260_t0,N4260_t1,N4260_t2,N4266_t0,N4266_t1,
     N957_t0,N957_t1,N4269_t0,N4269_t1,N4269_t2,N4278_t0,N4278_t1,N4275_t0,N4275_t1,N4281_t0,
     N4281_t1,N4281_t2,N4287_t0,N4287_t1,N1200_t0,N1200_t1,N4290_t0,N4290_t1,N4290_t2,N4294_t0,
     N4294_t1,N4294_t2,N4298_t0,N4298_t1,N4298_t2,N4302_t0,N4302_t1,N4302_t2,N4306_t0,N4306_t1,
     N4306_t2,N4310_t0,N4310_t1,N4310_t2,N4314_t0,N4314_t1,N4314_t2,N4320_t0,N4320_t1,N909_t0,
     N909_t1,N4323_t0,N4323_t1,N4323_t2,N4332_t0,N4332_t1,N4329_t0,N4329_t1,N4335_t0,N4335_t1,
     N4335_t2,N4341_t0,N4341_t1,N1152_t0,N1152_t1,N4344_t0,N4344_t1,N4344_t2,N1296_t0,N1296_t1,
     N4350_t0,N4350_t1,N4365_t0,N4365_t1,N861_t0,N861_t1,N4368_t0,N4368_t1,N4368_t2,N4377_t0,
     N4377_t1,N4374_t0,N4374_t1,N4380_t0,N4380_t1,N4380_t2,N4386_t0,N4386_t1,N1104_t0,N1104_t1,
     N4389_t0,N4389_t1,N4389_t2,N4398_t0,N4398_t1,N4395_t0,N4395_t1,N4401_t0,N4401_t1,N4401_t2,
     N4405_t0,N4405_t1,N573_t0,N573_t1,N4408_t0,N4408_t1,N621_t0,N621_t1,N4411_t0,N4411_t1,
     N669_t0,N669_t1,N4414_t0,N4414_t1,N717_t0,N717_t1,N4417_t0,N4417_t1,N765_t0,N765_t1,
     N4420_t0,N4420_t1,N813_t0,N813_t1,N4423_t0,N4423_t1,N4423_t2,N4432_t0,N4432_t1,N4429_t0,
     N4429_t1,N4435_t0,N4435_t1,N4435_t2,N4441_t0,N4441_t1,N1056_t0,N1056_t1,N4444_t0,N4444_t1,
     N4444_t2,N4453_t0,N4453_t1,N4450_t0,N4450_t1,N4456_t0,N4456_t1,N4456_t2,N4462_t0,N4462_t1,
     N4462_t2,N4466_t0,N4466_t1,N4466_t2,N4470_t0,N4470_t1,N4470_t2,N4474_t0,N4474_t1,N4474_t2,
     N4478_t0,N4478_t1,N4478_t2,N4482_t0,N4482_t1,N4482_t2,N4491_t0,N4491_t1,N4488_t0,N4488_t1,
     N4494_t0,N4494_t1,N4494_t2,N4500_t0,N4500_t1,N1008_t0,N1008_t1,N4503_t0,N4503_t1,N4503_t2,
     N4512_t0,N4512_t1,N4509_t0,N4509_t1,N4515_t0,N4515_t1,N4515_t2,N4521_t0,N4521_t1,N1251_t0,
     N1251_t1,N4554_t0,N4554_t1,N4551_t0,N4551_t1,N4557_t0,N4557_t1,N4557_t2,N4563_t0,N4563_t1,
     N960_t0,N960_t1,N4566_t0,N4566_t1,N4566_t2,N4575_t0,N4575_t1,N4572_t0,N4572_t1,N4578_t0,
     N4578_t1,N4578_t2,N4584_t0,N4584_t1,N1203_t0,N1203_t1,N4587_t0,N4587_t1,N4587_t2,N4592_t0,
     N4592_t1,N4526_t0,N4526_t1,N4595_t0,N4595_t1,N4531_t0,N4531_t1,N4598_t0,N4598_t1,N4536_t0,
     N4536_t1,N4601_t0,N4601_t1,N4541_t0,N4541_t1,N4604_t0,N4604_t1,N4546_t0,N4546_t1,N4607_t0,
     N4607_t1,N4607_t2,N4613_t0,N4613_t1,N912_t0,N912_t1,N4616_t0,N4616_t1,N4616_t2,N4625_t0,
     N4625_t1,N4622_t0,N4622_t1,N4628_t0,N4628_t1,N4628_t2,N4634_t0,N4634_t1,N1155_t0,N1155_t1,
     N4637_t0,N4637_t1,N4637_t2,N1299_t0,N1299_t1,N4643_t0,N4643_t1,N4646_t0,N4646_t1,N4646_t2,
     N4650_t0,N4650_t1,N4650_t2,N4654_t0,N4654_t1,N4654_t2,N4658_t0,N4658_t1,N4658_t2,N4662_t0,
     N4662_t1,N4662_t2,N4668_t0,N4668_t1,N864_t0,N864_t1,N4671_t0,N4671_t1,N4671_t2,N4680_t0,
     N4680_t1,N4677_t0,N4677_t1,N4683_t0,N4683_t1,N4683_t2,N4689_t0,N4689_t1,N1107_t0,N1107_t1,
     N4692_t0,N4692_t1,N4692_t2,N4701_t0,N4701_t1,N4698_t0,N4698_t1,N4704_t0,N4704_t1,N4704_t2,
     N4718_t0,N4718_t1,N816_t0,N816_t1,N4721_t0,N4721_t1,N4721_t2,N4730_t0,N4730_t1,N4727_t0,
     N4727_t1,N4733_t0,N4733_t1,N4733_t2,N4739_t0,N4739_t1,N1059_t0,N1059_t1,N4742_t0,N4742_t1,
     N4742_t2,N4751_t0,N4751_t1,N4748_t0,N4748_t1,N4754_t0,N4754_t1,N4754_t2,N4760_t0,N4760_t1,
     N576_t0,N576_t1,N4763_t0,N4763_t1,N624_t0,N624_t1,N4766_t0,N4766_t1,N672_t0,N672_t1,
     N4769_t0,N4769_t1,N720_t0,N720_t1,N4772_t0,N4772_t1,N768_t0,N768_t1,N4775_t0,N4775_t1,
     N4775_t2,N4784_t0,N4784_t1,N4781_t0,N4781_t1,N4787_t0,N4787_t1,N4787_t2,N4793_t0,N4793_t1,
     N1011_t0,N1011_t1,N4796_t0,N4796_t1,N4796_t2,N4805_t0,N4805_t1,N4802_t0,N4802_t1,N4808_t0,
     N4808_t1,N4808_t2,N4814_t0,N4814_t1,N1254_t0,N1254_t1,N4817_t0,N4817_t1,N4817_t2,N4821_t0,
     N4821_t1,N4821_t2,N4825_t0,N4825_t1,N4825_t2,N4829_t0,N4829_t1,N4829_t2,N4833_t0,N4833_t1,
     N4833_t2,N4842_t0,N4842_t1,N4839_t0,N4839_t1,N4845_t0,N4845_t1,N4845_t2,N4851_t0,N4851_t1,
     N963_t0,N963_t1,N4854_t0,N4854_t1,N4854_t2,N4863_t0,N4863_t1,N4860_t0,N4860_t1,N4866_t0,
     N4866_t1,N4866_t2,N4872_t0,N4872_t1,N1206_t0,N1206_t1,N4875_t0,N4875_t1,N4875_t2,N4904_t0,
     N4904_t1,N4901_t0,N4901_t1,N4907_t0,N4907_t1,N4907_t2,N4913_t0,N4913_t1,N915_t0,N915_t1,
     N4916_t0,N4916_t1,N4916_t2,N4925_t0,N4925_t1,N4922_t0,N4922_t1,N4928_t0,N4928_t1,N4928_t2,
     N4934_t0,N4934_t1,N1158_t0,N1158_t1,N4937_t0,N4937_t1,N4937_t2,N1302_t0,N1302_t1,N4943_t0,
     N4943_t1,N4947_t0,N4947_t1,N4881_t0,N4881_t1,N4950_t0,N4950_t1,N4886_t0,N4886_t1,N4953_t0,
     N4953_t1,N4891_t0,N4891_t1,N4956_t0,N4956_t1,N4896_t0,N4896_t1,N4959_t0,N4959_t1,N4959_t2,
     N4965_t0,N4965_t1,N867_t0,N867_t1,N4968_t0,N4968_t1,N4968_t2,N4977_t0,N4977_t1,N4974_t0,
     N4974_t1,N4980_t0,N4980_t1,N4980_t2,N4986_t0,N4986_t1,N1110_t0,N1110_t1,N4989_t0,N4989_t1,
     N4989_t2,N4998_t0,N4998_t1,N4995_t0,N4995_t1,N5001_t0,N5001_t1,N5001_t2,N5005_t0,N5005_t1,
     N5005_t2,N5009_t0,N5009_t1,N5009_t2,N5013_t0,N5013_t1,N5013_t2,N5017_t0,N5017_t1,N5017_t2,
     N5023_t0,N5023_t1,N819_t0,N819_t1,N5026_t0,N5026_t1,N5026_t2,N5035_t0,N5035_t1,N5032_t0,
     N5032_t1,N5038_t0,N5038_t1,N5038_t2,N5044_t0,N5044_t1,N1062_t0,N1062_t1,N5047_t0,N5047_t1,
     N5047_t2,N5056_t0,N5056_t1,N5053_t0,N5053_t1,N5059_t0,N5059_t1,N5059_t2,N5073_t0,N5073_t1,
     N771_t0,N771_t1,N5076_t0,N5076_t1,N5076_t2,N5085_t0,N5085_t1,N5082_t0,N5082_t1,N5088_t0,
     N5088_t1,N5088_t2,N5094_t0,N5094_t1,N1014_t0,N1014_t1,N5097_t0,N5097_t1,N5097_t2,N5106_t0,
     N5106_t1,N5103_t0,N5103_t1,N5109_t0,N5109_t1,N5109_t2,N5115_t0,N5115_t1,N1257_t0,N1257_t1,
     N5118_t0,N5118_t1,N579_t0,N579_t1,N5121_t0,N5121_t1,N627_t0,N627_t1,N5124_t0,N5124_t1,
     N675_t0,N675_t1,N5127_t0,N5127_t1,N723_t0,N723_t1,N5130_t0,N5130_t1,N5130_t2,N5139_t0,
     N5139_t1,N5136_t0,N5136_t1,N5142_t0,N5142_t1,N5142_t2,N5148_t0,N5148_t1,N966_t0,N966_t1,
     N5151_t0,N5151_t1,N5151_t2,N5160_t0,N5160_t1,N5157_t0,N5157_t1,N5163_t0,N5163_t1,N5163_t2,
     N5169_t0,N5169_t1,N1209_t0,N1209_t1,N5172_t0,N5172_t1,N5172_t2,N5176_t0,N5176_t1,N5176_t2,
     N5180_t0,N5180_t1,N5180_t2,N5184_t0,N5184_t1,N5184_t2,N5188_t0,N5188_t1,N5188_t2,N5197_t0,
     N5197_t1,N5194_t0,N5194_t1,N5200_t0,N5200_t1,N5200_t2,N5206_t0,N5206_t1,N918_t0,N918_t1,
     N5209_t0,N5209_t1,N5209_t2,N5218_t0,N5218_t1,N5215_t0,N5215_t1,N5221_t0,N5221_t1,N5221_t2,
     N5227_t0,N5227_t1,N1161_t0,N1161_t1,N5230_t0,N5230_t1,N5230_t2,N1305_t0,N1305_t1,N5236_t0,
     N5236_t1,N5259_t0,N5259_t1,N5256_t0,N5256_t1,N5262_t0,N5262_t1,N5262_t2,N5268_t0,N5268_t1,
     N870_t0,N870_t1,N5271_t0,N5271_t1,N5271_t2,N5280_t0,N5280_t1,N5277_t0,N5277_t1,N5283_t0,
     N5283_t1,N5283_t2,N5289_t0,N5289_t1,N1113_t0,N1113_t1,N5292_t0,N5292_t1,N5292_t2,N5301_t0,
     N5301_t1,N5298_t0,N5298_t1,N5304_t0,N5304_t1,N5304_t2,N5309_t0,N5309_t1,N5241_t0,N5241_t1,
     N5312_t0,N5312_t1,N5246_t0,N5246_t1,N5315_t0,N5315_t1,N5251_t0,N5251_t1,N5318_t0,N5318_t1,
     N5318_t2,N5324_t0,N5324_t1,N822_t0,N822_t1,N5327_t0,N5327_t1,N5327_t2,N5336_t0,N5336_t1,
     N5333_t0,N5333_t1,N5339_t0,N5339_t1,N5339_t2,N5345_t0,N5345_t1,N1065_t0,N1065_t1,N5348_t0,
     N5348_t1,N5348_t2,N5357_t0,N5357_t1,N5354_t0,N5354_t1,N5360_t0,N5360_t1,N5360_t2,N5366_t0,
     N5366_t1,N5366_t2,N5370_t0,N5370_t1,N5370_t2,N5374_t0,N5374_t1,N5374_t2,N5380_t0,N5380_t1,
     N774_t0,N774_t1,N5383_t0,N5383_t1,N5383_t2,N5392_t0,N5392_t1,N5389_t0,N5389_t1,N5395_t0,
     N5395_t1,N5395_t2,N5401_t0,N5401_t1,N1017_t0,N1017_t1,N5404_t0,N5404_t1,N5404_t2,N5413_t0,
     N5413_t1,N5410_t0,N5410_t1,N5416_t0,N5416_t1,N5416_t2,N5422_t0,N5422_t1,N1260_t0,N1260_t1,
     N5431_t0,N5431_t1,N726_t0,N726_t1,N5434_t0,N5434_t1,N5434_t2,N5443_t0,N5443_t1,N5440_t0,
     N5440_t1,N5446_t0,N5446_t1,N5446_t2,N5452_t0,N5452_t1,N969_t0,N969_t1,N5455_t0,N5455_t1,
     N5455_t2,N5464_t0,N5464_t1,N5461_t0,N5461_t1,N5467_t0,N5467_t1,N5467_t2,N5473_t0,N5473_t1,
     N1212_t0,N1212_t1,N5476_t0,N5476_t1,N5476_t2,N5480_t0,N5480_t1,N582_t0,N582_t1,N5483_t0,
     N5483_t1,N630_t0,N630_t1,N5486_t0,N5486_t1,N678_t0,N678_t1,N5489_t0,N5489_t1,N5489_t2,
     N5498_t0,N5498_t1,N5495_t0,N5495_t1,N5501_t0,N5501_t1,N5501_t2,N5507_t0,N5507_t1,N921_t0,
     N921_t1,N5510_t0,N5510_t1,N5510_t2,N5519_t0,N5519_t1,N5516_t0,N5516_t1,N5522_t0,N5522_t1,
     N5522_t2,N5528_t0,N5528_t1,N1164_t0,N1164_t1,N5531_t0,N5531_t1,N5531_t2,N1308_t0,N1308_t1,
     N5537_t0,N5537_t1,N5540_t0,N5540_t1,N5540_t2,N5544_t0,N5544_t1,N5544_t2,N5548_t0,N5548_t1,
     N5548_t2,N5557_t0,N5557_t1,N5554_t0,N5554_t1,N5560_t0,N5560_t1,N5560_t2,N5566_t0,N5566_t1,
     N873_t0,N873_t1,N5569_t0,N5569_t1,N5569_t2,N5578_t0,N5578_t1,N5575_t0,N5575_t1,N5581_t0,
     N5581_t1,N5581_t2,N5587_t0,N5587_t1,N1116_t0,N1116_t1,N5590_t0,N5590_t1,N5590_t2,N5599_t0,
     N5599_t1,N5596_t0,N5596_t1,N5602_t0,N5602_t1,N5602_t2,N5621_t0,N5621_t1,N5618_t0,N5618_t1,
     N5624_t0,N5624_t1,N5624_t2,N5630_t0,N5630_t1,N825_t0,N825_t1,N5633_t0,N5633_t1,N5633_t2,
     N5642_t0,N5642_t1,N5639_t0,N5639_t1,N5645_t0,N5645_t1,N5645_t2,N5651_t0,N5651_t1,N1068_t0,
     N1068_t1,N5654_t0,N5654_t1,N5654_t2,N5663_t0,N5663_t1,N5660_t0,N5660_t1,N5666_t0,N5666_t1,
     N5666_t2,N5673_t0,N5673_t1,N5608_t0,N5608_t1,N5676_t0,N5676_t1,N5613_t0,N5613_t1,N5679_t0,
     N5679_t1,N5679_t2,N5685_t0,N5685_t1,N777_t0,N777_t1,N5688_t0,N5688_t1,N5688_t2,N5697_t0,
     N5697_t1,N5694_t0,N5694_t1,N5700_t0,N5700_t1,N5700_t2,N5706_t0,N5706_t1,N1020_t0,N1020_t1,
     N5709_t0,N5709_t1,N5709_t2,N5718_t0,N5718_t1,N5715_t0,N5715_t1,N5721_t0,N5721_t1,N5721_t2,
     N5730_t0,N5730_t1,N5730_t2,N5734_t0,N5734_t1,N5734_t2,N5740_t0,N5740_t1,N729_t0,N729_t1,
     N5743_t0,N5743_t1,N5743_t2,N5752_t0,N5752_t1,N5749_t0,N5749_t1,N5755_t0,N5755_t1,N5755_t2,
     N5761_t0,N5761_t1,N972_t0,N972_t1,N5764_t0,N5764_t1,N5764_t2,N5773_t0,N5773_t1,N5770_t0,
     N5770_t1,N5776_t0,N5776_t1,N5776_t2,N5789_t0,N5789_t1,N681_t0,N681_t1,N5792_t0,N5792_t1,
     N5792_t2,N5801_t0,N5801_t1,N5798_t0,N5798_t1,N5804_t0,N5804_t1,N5804_t2,N5810_t0,N5810_t1,
     N924_t0,N924_t1,N5813_t0,N5813_t1,N5813_t2,N5822_t0,N5822_t1,N5819_t0,N5819_t1,N5825_t0,
     N5825_t1,N5825_t2,N5834_t0,N5834_t1,N585_t0,N585_t1,N5837_t0,N5837_t1,N633_t0,N633_t1,
     N5840_t0,N5840_t1,N5840_t2,N5849_t0,N5849_t1,N5846_t0,N5846_t1,N5852_t0,N5852_t1,N5852_t2,
     N5858_t0,N5858_t1,N876_t0,N876_t1,N5861_t0,N5861_t1,N5861_t2,N5870_t0,N5870_t1,N5867_t0,
     N5867_t1,N5873_t0,N5873_t1,N5873_t2,N5882_t0,N5882_t1,N5882_t2,N5886_t0,N5886_t1,N5886_t2,
     N5895_t0,N5895_t1,N5892_t0,N5892_t1,N5898_t0,N5898_t1,N5898_t2,N5904_t0,N5904_t1,N828_t0,
     N828_t1,N5907_t0,N5907_t1,N5907_t2,N5916_t0,N5916_t1,N5913_t0,N5913_t1,N5919_t0,N5919_t1,
     N5919_t2,N5938_t0,N5938_t1,N5935_t0,N5935_t1,N5941_t0,N5941_t1,N5941_t2,N5947_t0,N5947_t1,
     N780_t0,N780_t1,N5950_t0,N5950_t1,N5950_t2,N5959_t0,N5959_t1,N5956_t0,N5956_t1,N5962_t0,
     N5962_t1,N5962_t2,N5972_t0,N5972_t1,N5930_t0,N5930_t1,N5975_t0,N5975_t1,N5975_t2,N5981_t0,
     N5981_t1,N732_t0,N732_t1,N5984_t0,N5984_t1,N5984_t2,N5993_t0,N5993_t1,N5990_t0,N5990_t1,
     N5996_t0,N5996_t1,N5996_t2,N6005_t0,N6005_t1,N6005_t2,N6011_t0,N6011_t1,N684_t0,N684_t1,
     N6014_t0,N6014_t1,N6014_t2,N6023_t0,N6023_t1,N6020_t0,N6020_t1,N6026_t0,N6026_t1,N6026_t2,
     N6037_t0,N6037_t1,N636_t0,N636_t1,N6040_t0,N6040_t1,N6040_t2,N6049_t0,N6049_t1,N6046_t0,
     N6046_t1,N6052_t0,N6052_t1,N6052_t2,N6061_t0,N6061_t1,N588_t0,N588_t1,N6064_t0,N6064_t1,
     N6064_t2,N6073_t0,N6073_t1,N6070_t0,N6070_t1,N6076_t0,N6076_t1,N6076_t2,N6085_t0,N6085_t1,
     N6085_t2,N6094_t0,N6094_t1,N6091_t0,N6091_t1,N6097_t0,N6097_t1,N6097_t2,N6111_t0,N6111_t1,
     N6108_t0,N6108_t1,N6114_t0,N6114_t1,N6114_t2,N6124_t0,N6124_t1,N6124_t2,N6138_t0,N6138_t1,
     N6141_t0,N6141_t1,N6141_t2,N6135_t0,N6135_t1,N6147_t0,N6147_t1,N6151_t0,N6151_t1,N6151_t2,
     N6130_t0,N6130_t1,N6157_t0,N6157_t1,N6161_t0,N6161_t1,N6161_t2,N6120_t0,N6120_t1,N6167_t0,
     N6167_t1,N6171_t0,N6171_t1,N6171_t2,N6103_t0,N6103_t1,N6177_t0,N6177_t1,N6181_t0,N6181_t1,
     N6181_t2,N6082_t0,N6082_t1,N6187_t0,N6187_t1,N6191_t0,N6191_t1,N6191_t2,N6058_t0,N6058_t1,
     N6197_t0,N6197_t1,N6201_t0,N6201_t1,N6201_t2,N6032_t0,N6032_t1,N6207_t0,N6207_t1,N6211_t0,
     N6211_t1,N6211_t2,N6002_t0,N6002_t1,N6217_t0,N6217_t1,N6221_t0,N6221_t1,N6221_t2,N5968_t0,
     N5968_t1,N6227_t0,N6227_t1,N6231_t0,N6231_t1,N6231_t2,N5925_t0,N5925_t1,N6237_t0,N6237_t1,
     N6241_t0,N6241_t1,N6241_t2,N5879_t0,N5879_t1,N6247_t0,N6247_t1,N6251_t0,N6251_t1,N6251_t2,
     N5831_t0,N5831_t1,N6257_t0,N6257_t1,N6261_t0,N6261_t1,N6261_t2,N5782_t0,N5782_t1,N6267_t0,
     N6267_t1,N6271_t0,N6271_t1,N6271_t2,N5727_t0,N5727_t1,N6277_t0,N6277_t1,N6281_t0,N6281_t1,
     N6281_t2;
reg [3839:0] FEN;
fim FAN_N1_0 ( .fault(fault), .net(N1), .FEN(FEN[0]), .op(N1_t0) );
fim FAN_N1_1 ( .fault(fault), .net(N1), .FEN(FEN[1]), .op(N1_t1) );
fim FAN_N1_2 ( .fault(fault), .net(N1), .FEN(FEN[2]), .op(N1_t2) );
fim FAN_N1_3 ( .fault(fault), .net(N1), .FEN(FEN[3]), .op(N1_t3) );
fim FAN_N1_4 ( .fault(fault), .net(N1), .FEN(FEN[4]), .op(N1_t4) );
fim FAN_N1_5 ( .fault(fault), .net(N1), .FEN(FEN[5]), .op(N1_t5) );
fim FAN_N1_6 ( .fault(fault), .net(N1), .FEN(FEN[6]), .op(N1_t6) );
fim FAN_N1_7 ( .fault(fault), .net(N1), .FEN(FEN[7]), .op(N1_t7) );
fim FAN_N1_8 ( .fault(fault), .net(N1), .FEN(FEN[8]), .op(N1_t8) );
fim FAN_N1_9 ( .fault(fault), .net(N1), .FEN(FEN[9]), .op(N1_t9) );
fim FAN_N1_10 ( .fault(fault), .net(N1), .FEN(FEN[10]), .op(N1_t10) );
fim FAN_N1_11 ( .fault(fault), .net(N1), .FEN(FEN[11]), .op(N1_t11) );
fim FAN_N1_12 ( .fault(fault), .net(N1), .FEN(FEN[12]), .op(N1_t12) );
fim FAN_N1_13 ( .fault(fault), .net(N1), .FEN(FEN[13]), .op(N1_t13) );
fim FAN_N1_14 ( .fault(fault), .net(N1), .FEN(FEN[14]), .op(N1_t14) );
fim FAN_N1_15 ( .fault(fault), .net(N1), .FEN(FEN[15]), .op(N1_t15) );
fim FAN_N273_0 ( .fault(fault), .net(N273), .FEN(FEN[16]), .op(N273_t0) );
fim FAN_N273_1 ( .fault(fault), .net(N273), .FEN(FEN[17]), .op(N273_t1) );
fim FAN_N273_2 ( .fault(fault), .net(N273), .FEN(FEN[18]), .op(N273_t2) );
fim FAN_N273_3 ( .fault(fault), .net(N273), .FEN(FEN[19]), .op(N273_t3) );
fim FAN_N273_4 ( .fault(fault), .net(N273), .FEN(FEN[20]), .op(N273_t4) );
fim FAN_N273_5 ( .fault(fault), .net(N273), .FEN(FEN[21]), .op(N273_t5) );
fim FAN_N273_6 ( .fault(fault), .net(N273), .FEN(FEN[22]), .op(N273_t6) );
fim FAN_N273_7 ( .fault(fault), .net(N273), .FEN(FEN[23]), .op(N273_t7) );
fim FAN_N273_8 ( .fault(fault), .net(N273), .FEN(FEN[24]), .op(N273_t8) );
fim FAN_N273_9 ( .fault(fault), .net(N273), .FEN(FEN[25]), .op(N273_t9) );
fim FAN_N273_10 ( .fault(fault), .net(N273), .FEN(FEN[26]), .op(N273_t10) );
fim FAN_N273_11 ( .fault(fault), .net(N273), .FEN(FEN[27]), .op(N273_t11) );
fim FAN_N273_12 ( .fault(fault), .net(N273), .FEN(FEN[28]), .op(N273_t12) );
fim FAN_N273_13 ( .fault(fault), .net(N273), .FEN(FEN[29]), .op(N273_t13) );
fim FAN_N273_14 ( .fault(fault), .net(N273), .FEN(FEN[30]), .op(N273_t14) );
fim FAN_N273_15 ( .fault(fault), .net(N273), .FEN(FEN[31]), .op(N273_t15) );
fim FAN_N290_0 ( .fault(fault), .net(N290), .FEN(FEN[32]), .op(N290_t0) );
fim FAN_N290_1 ( .fault(fault), .net(N290), .FEN(FEN[33]), .op(N290_t1) );
fim FAN_N290_2 ( .fault(fault), .net(N290), .FEN(FEN[34]), .op(N290_t2) );
fim FAN_N290_3 ( .fault(fault), .net(N290), .FEN(FEN[35]), .op(N290_t3) );
fim FAN_N290_4 ( .fault(fault), .net(N290), .FEN(FEN[36]), .op(N290_t4) );
fim FAN_N290_5 ( .fault(fault), .net(N290), .FEN(FEN[37]), .op(N290_t5) );
fim FAN_N290_6 ( .fault(fault), .net(N290), .FEN(FEN[38]), .op(N290_t6) );
fim FAN_N290_7 ( .fault(fault), .net(N290), .FEN(FEN[39]), .op(N290_t7) );
fim FAN_N290_8 ( .fault(fault), .net(N290), .FEN(FEN[40]), .op(N290_t8) );
fim FAN_N290_9 ( .fault(fault), .net(N290), .FEN(FEN[41]), .op(N290_t9) );
fim FAN_N290_10 ( .fault(fault), .net(N290), .FEN(FEN[42]), .op(N290_t10) );
fim FAN_N290_11 ( .fault(fault), .net(N290), .FEN(FEN[43]), .op(N290_t11) );
fim FAN_N290_12 ( .fault(fault), .net(N290), .FEN(FEN[44]), .op(N290_t12) );
fim FAN_N290_13 ( .fault(fault), .net(N290), .FEN(FEN[45]), .op(N290_t13) );
fim FAN_N290_14 ( .fault(fault), .net(N290), .FEN(FEN[46]), .op(N290_t14) );
fim FAN_N290_15 ( .fault(fault), .net(N290), .FEN(FEN[47]), .op(N290_t15) );
fim FAN_N307_0 ( .fault(fault), .net(N307), .FEN(FEN[48]), .op(N307_t0) );
fim FAN_N307_1 ( .fault(fault), .net(N307), .FEN(FEN[49]), .op(N307_t1) );
fim FAN_N307_2 ( .fault(fault), .net(N307), .FEN(FEN[50]), .op(N307_t2) );
fim FAN_N307_3 ( .fault(fault), .net(N307), .FEN(FEN[51]), .op(N307_t3) );
fim FAN_N307_4 ( .fault(fault), .net(N307), .FEN(FEN[52]), .op(N307_t4) );
fim FAN_N307_5 ( .fault(fault), .net(N307), .FEN(FEN[53]), .op(N307_t5) );
fim FAN_N307_6 ( .fault(fault), .net(N307), .FEN(FEN[54]), .op(N307_t6) );
fim FAN_N307_7 ( .fault(fault), .net(N307), .FEN(FEN[55]), .op(N307_t7) );
fim FAN_N307_8 ( .fault(fault), .net(N307), .FEN(FEN[56]), .op(N307_t8) );
fim FAN_N307_9 ( .fault(fault), .net(N307), .FEN(FEN[57]), .op(N307_t9) );
fim FAN_N307_10 ( .fault(fault), .net(N307), .FEN(FEN[58]), .op(N307_t10) );
fim FAN_N307_11 ( .fault(fault), .net(N307), .FEN(FEN[59]), .op(N307_t11) );
fim FAN_N307_12 ( .fault(fault), .net(N307), .FEN(FEN[60]), .op(N307_t12) );
fim FAN_N307_13 ( .fault(fault), .net(N307), .FEN(FEN[61]), .op(N307_t13) );
fim FAN_N307_14 ( .fault(fault), .net(N307), .FEN(FEN[62]), .op(N307_t14) );
fim FAN_N307_15 ( .fault(fault), .net(N307), .FEN(FEN[63]), .op(N307_t15) );
fim FAN_N324_0 ( .fault(fault), .net(N324), .FEN(FEN[64]), .op(N324_t0) );
fim FAN_N324_1 ( .fault(fault), .net(N324), .FEN(FEN[65]), .op(N324_t1) );
fim FAN_N324_2 ( .fault(fault), .net(N324), .FEN(FEN[66]), .op(N324_t2) );
fim FAN_N324_3 ( .fault(fault), .net(N324), .FEN(FEN[67]), .op(N324_t3) );
fim FAN_N324_4 ( .fault(fault), .net(N324), .FEN(FEN[68]), .op(N324_t4) );
fim FAN_N324_5 ( .fault(fault), .net(N324), .FEN(FEN[69]), .op(N324_t5) );
fim FAN_N324_6 ( .fault(fault), .net(N324), .FEN(FEN[70]), .op(N324_t6) );
fim FAN_N324_7 ( .fault(fault), .net(N324), .FEN(FEN[71]), .op(N324_t7) );
fim FAN_N324_8 ( .fault(fault), .net(N324), .FEN(FEN[72]), .op(N324_t8) );
fim FAN_N324_9 ( .fault(fault), .net(N324), .FEN(FEN[73]), .op(N324_t9) );
fim FAN_N324_10 ( .fault(fault), .net(N324), .FEN(FEN[74]), .op(N324_t10) );
fim FAN_N324_11 ( .fault(fault), .net(N324), .FEN(FEN[75]), .op(N324_t11) );
fim FAN_N324_12 ( .fault(fault), .net(N324), .FEN(FEN[76]), .op(N324_t12) );
fim FAN_N324_13 ( .fault(fault), .net(N324), .FEN(FEN[77]), .op(N324_t13) );
fim FAN_N324_14 ( .fault(fault), .net(N324), .FEN(FEN[78]), .op(N324_t14) );
fim FAN_N324_15 ( .fault(fault), .net(N324), .FEN(FEN[79]), .op(N324_t15) );
fim FAN_N341_0 ( .fault(fault), .net(N341), .FEN(FEN[80]), .op(N341_t0) );
fim FAN_N341_1 ( .fault(fault), .net(N341), .FEN(FEN[81]), .op(N341_t1) );
fim FAN_N341_2 ( .fault(fault), .net(N341), .FEN(FEN[82]), .op(N341_t2) );
fim FAN_N341_3 ( .fault(fault), .net(N341), .FEN(FEN[83]), .op(N341_t3) );
fim FAN_N341_4 ( .fault(fault), .net(N341), .FEN(FEN[84]), .op(N341_t4) );
fim FAN_N341_5 ( .fault(fault), .net(N341), .FEN(FEN[85]), .op(N341_t5) );
fim FAN_N341_6 ( .fault(fault), .net(N341), .FEN(FEN[86]), .op(N341_t6) );
fim FAN_N341_7 ( .fault(fault), .net(N341), .FEN(FEN[87]), .op(N341_t7) );
fim FAN_N341_8 ( .fault(fault), .net(N341), .FEN(FEN[88]), .op(N341_t8) );
fim FAN_N341_9 ( .fault(fault), .net(N341), .FEN(FEN[89]), .op(N341_t9) );
fim FAN_N341_10 ( .fault(fault), .net(N341), .FEN(FEN[90]), .op(N341_t10) );
fim FAN_N341_11 ( .fault(fault), .net(N341), .FEN(FEN[91]), .op(N341_t11) );
fim FAN_N341_12 ( .fault(fault), .net(N341), .FEN(FEN[92]), .op(N341_t12) );
fim FAN_N341_13 ( .fault(fault), .net(N341), .FEN(FEN[93]), .op(N341_t13) );
fim FAN_N341_14 ( .fault(fault), .net(N341), .FEN(FEN[94]), .op(N341_t14) );
fim FAN_N341_15 ( .fault(fault), .net(N341), .FEN(FEN[95]), .op(N341_t15) );
fim FAN_N358_0 ( .fault(fault), .net(N358), .FEN(FEN[96]), .op(N358_t0) );
fim FAN_N358_1 ( .fault(fault), .net(N358), .FEN(FEN[97]), .op(N358_t1) );
fim FAN_N358_2 ( .fault(fault), .net(N358), .FEN(FEN[98]), .op(N358_t2) );
fim FAN_N358_3 ( .fault(fault), .net(N358), .FEN(FEN[99]), .op(N358_t3) );
fim FAN_N358_4 ( .fault(fault), .net(N358), .FEN(FEN[100]), .op(N358_t4) );
fim FAN_N358_5 ( .fault(fault), .net(N358), .FEN(FEN[101]), .op(N358_t5) );
fim FAN_N358_6 ( .fault(fault), .net(N358), .FEN(FEN[102]), .op(N358_t6) );
fim FAN_N358_7 ( .fault(fault), .net(N358), .FEN(FEN[103]), .op(N358_t7) );
fim FAN_N358_8 ( .fault(fault), .net(N358), .FEN(FEN[104]), .op(N358_t8) );
fim FAN_N358_9 ( .fault(fault), .net(N358), .FEN(FEN[105]), .op(N358_t9) );
fim FAN_N358_10 ( .fault(fault), .net(N358), .FEN(FEN[106]), .op(N358_t10) );
fim FAN_N358_11 ( .fault(fault), .net(N358), .FEN(FEN[107]), .op(N358_t11) );
fim FAN_N358_12 ( .fault(fault), .net(N358), .FEN(FEN[108]), .op(N358_t12) );
fim FAN_N358_13 ( .fault(fault), .net(N358), .FEN(FEN[109]), .op(N358_t13) );
fim FAN_N358_14 ( .fault(fault), .net(N358), .FEN(FEN[110]), .op(N358_t14) );
fim FAN_N358_15 ( .fault(fault), .net(N358), .FEN(FEN[111]), .op(N358_t15) );
fim FAN_N375_0 ( .fault(fault), .net(N375), .FEN(FEN[112]), .op(N375_t0) );
fim FAN_N375_1 ( .fault(fault), .net(N375), .FEN(FEN[113]), .op(N375_t1) );
fim FAN_N375_2 ( .fault(fault), .net(N375), .FEN(FEN[114]), .op(N375_t2) );
fim FAN_N375_3 ( .fault(fault), .net(N375), .FEN(FEN[115]), .op(N375_t3) );
fim FAN_N375_4 ( .fault(fault), .net(N375), .FEN(FEN[116]), .op(N375_t4) );
fim FAN_N375_5 ( .fault(fault), .net(N375), .FEN(FEN[117]), .op(N375_t5) );
fim FAN_N375_6 ( .fault(fault), .net(N375), .FEN(FEN[118]), .op(N375_t6) );
fim FAN_N375_7 ( .fault(fault), .net(N375), .FEN(FEN[119]), .op(N375_t7) );
fim FAN_N375_8 ( .fault(fault), .net(N375), .FEN(FEN[120]), .op(N375_t8) );
fim FAN_N375_9 ( .fault(fault), .net(N375), .FEN(FEN[121]), .op(N375_t9) );
fim FAN_N375_10 ( .fault(fault), .net(N375), .FEN(FEN[122]), .op(N375_t10) );
fim FAN_N375_11 ( .fault(fault), .net(N375), .FEN(FEN[123]), .op(N375_t11) );
fim FAN_N375_12 ( .fault(fault), .net(N375), .FEN(FEN[124]), .op(N375_t12) );
fim FAN_N375_13 ( .fault(fault), .net(N375), .FEN(FEN[125]), .op(N375_t13) );
fim FAN_N375_14 ( .fault(fault), .net(N375), .FEN(FEN[126]), .op(N375_t14) );
fim FAN_N375_15 ( .fault(fault), .net(N375), .FEN(FEN[127]), .op(N375_t15) );
fim FAN_N392_0 ( .fault(fault), .net(N392), .FEN(FEN[128]), .op(N392_t0) );
fim FAN_N392_1 ( .fault(fault), .net(N392), .FEN(FEN[129]), .op(N392_t1) );
fim FAN_N392_2 ( .fault(fault), .net(N392), .FEN(FEN[130]), .op(N392_t2) );
fim FAN_N392_3 ( .fault(fault), .net(N392), .FEN(FEN[131]), .op(N392_t3) );
fim FAN_N392_4 ( .fault(fault), .net(N392), .FEN(FEN[132]), .op(N392_t4) );
fim FAN_N392_5 ( .fault(fault), .net(N392), .FEN(FEN[133]), .op(N392_t5) );
fim FAN_N392_6 ( .fault(fault), .net(N392), .FEN(FEN[134]), .op(N392_t6) );
fim FAN_N392_7 ( .fault(fault), .net(N392), .FEN(FEN[135]), .op(N392_t7) );
fim FAN_N392_8 ( .fault(fault), .net(N392), .FEN(FEN[136]), .op(N392_t8) );
fim FAN_N392_9 ( .fault(fault), .net(N392), .FEN(FEN[137]), .op(N392_t9) );
fim FAN_N392_10 ( .fault(fault), .net(N392), .FEN(FEN[138]), .op(N392_t10) );
fim FAN_N392_11 ( .fault(fault), .net(N392), .FEN(FEN[139]), .op(N392_t11) );
fim FAN_N392_12 ( .fault(fault), .net(N392), .FEN(FEN[140]), .op(N392_t12) );
fim FAN_N392_13 ( .fault(fault), .net(N392), .FEN(FEN[141]), .op(N392_t13) );
fim FAN_N392_14 ( .fault(fault), .net(N392), .FEN(FEN[142]), .op(N392_t14) );
fim FAN_N392_15 ( .fault(fault), .net(N392), .FEN(FEN[143]), .op(N392_t15) );
fim FAN_N409_0 ( .fault(fault), .net(N409), .FEN(FEN[144]), .op(N409_t0) );
fim FAN_N409_1 ( .fault(fault), .net(N409), .FEN(FEN[145]), .op(N409_t1) );
fim FAN_N409_2 ( .fault(fault), .net(N409), .FEN(FEN[146]), .op(N409_t2) );
fim FAN_N409_3 ( .fault(fault), .net(N409), .FEN(FEN[147]), .op(N409_t3) );
fim FAN_N409_4 ( .fault(fault), .net(N409), .FEN(FEN[148]), .op(N409_t4) );
fim FAN_N409_5 ( .fault(fault), .net(N409), .FEN(FEN[149]), .op(N409_t5) );
fim FAN_N409_6 ( .fault(fault), .net(N409), .FEN(FEN[150]), .op(N409_t6) );
fim FAN_N409_7 ( .fault(fault), .net(N409), .FEN(FEN[151]), .op(N409_t7) );
fim FAN_N409_8 ( .fault(fault), .net(N409), .FEN(FEN[152]), .op(N409_t8) );
fim FAN_N409_9 ( .fault(fault), .net(N409), .FEN(FEN[153]), .op(N409_t9) );
fim FAN_N409_10 ( .fault(fault), .net(N409), .FEN(FEN[154]), .op(N409_t10) );
fim FAN_N409_11 ( .fault(fault), .net(N409), .FEN(FEN[155]), .op(N409_t11) );
fim FAN_N409_12 ( .fault(fault), .net(N409), .FEN(FEN[156]), .op(N409_t12) );
fim FAN_N409_13 ( .fault(fault), .net(N409), .FEN(FEN[157]), .op(N409_t13) );
fim FAN_N409_14 ( .fault(fault), .net(N409), .FEN(FEN[158]), .op(N409_t14) );
fim FAN_N409_15 ( .fault(fault), .net(N409), .FEN(FEN[159]), .op(N409_t15) );
fim FAN_N426_0 ( .fault(fault), .net(N426), .FEN(FEN[160]), .op(N426_t0) );
fim FAN_N426_1 ( .fault(fault), .net(N426), .FEN(FEN[161]), .op(N426_t1) );
fim FAN_N426_2 ( .fault(fault), .net(N426), .FEN(FEN[162]), .op(N426_t2) );
fim FAN_N426_3 ( .fault(fault), .net(N426), .FEN(FEN[163]), .op(N426_t3) );
fim FAN_N426_4 ( .fault(fault), .net(N426), .FEN(FEN[164]), .op(N426_t4) );
fim FAN_N426_5 ( .fault(fault), .net(N426), .FEN(FEN[165]), .op(N426_t5) );
fim FAN_N426_6 ( .fault(fault), .net(N426), .FEN(FEN[166]), .op(N426_t6) );
fim FAN_N426_7 ( .fault(fault), .net(N426), .FEN(FEN[167]), .op(N426_t7) );
fim FAN_N426_8 ( .fault(fault), .net(N426), .FEN(FEN[168]), .op(N426_t8) );
fim FAN_N426_9 ( .fault(fault), .net(N426), .FEN(FEN[169]), .op(N426_t9) );
fim FAN_N426_10 ( .fault(fault), .net(N426), .FEN(FEN[170]), .op(N426_t10) );
fim FAN_N426_11 ( .fault(fault), .net(N426), .FEN(FEN[171]), .op(N426_t11) );
fim FAN_N426_12 ( .fault(fault), .net(N426), .FEN(FEN[172]), .op(N426_t12) );
fim FAN_N426_13 ( .fault(fault), .net(N426), .FEN(FEN[173]), .op(N426_t13) );
fim FAN_N426_14 ( .fault(fault), .net(N426), .FEN(FEN[174]), .op(N426_t14) );
fim FAN_N426_15 ( .fault(fault), .net(N426), .FEN(FEN[175]), .op(N426_t15) );
fim FAN_N443_0 ( .fault(fault), .net(N443), .FEN(FEN[176]), .op(N443_t0) );
fim FAN_N443_1 ( .fault(fault), .net(N443), .FEN(FEN[177]), .op(N443_t1) );
fim FAN_N443_2 ( .fault(fault), .net(N443), .FEN(FEN[178]), .op(N443_t2) );
fim FAN_N443_3 ( .fault(fault), .net(N443), .FEN(FEN[179]), .op(N443_t3) );
fim FAN_N443_4 ( .fault(fault), .net(N443), .FEN(FEN[180]), .op(N443_t4) );
fim FAN_N443_5 ( .fault(fault), .net(N443), .FEN(FEN[181]), .op(N443_t5) );
fim FAN_N443_6 ( .fault(fault), .net(N443), .FEN(FEN[182]), .op(N443_t6) );
fim FAN_N443_7 ( .fault(fault), .net(N443), .FEN(FEN[183]), .op(N443_t7) );
fim FAN_N443_8 ( .fault(fault), .net(N443), .FEN(FEN[184]), .op(N443_t8) );
fim FAN_N443_9 ( .fault(fault), .net(N443), .FEN(FEN[185]), .op(N443_t9) );
fim FAN_N443_10 ( .fault(fault), .net(N443), .FEN(FEN[186]), .op(N443_t10) );
fim FAN_N443_11 ( .fault(fault), .net(N443), .FEN(FEN[187]), .op(N443_t11) );
fim FAN_N443_12 ( .fault(fault), .net(N443), .FEN(FEN[188]), .op(N443_t12) );
fim FAN_N443_13 ( .fault(fault), .net(N443), .FEN(FEN[189]), .op(N443_t13) );
fim FAN_N443_14 ( .fault(fault), .net(N443), .FEN(FEN[190]), .op(N443_t14) );
fim FAN_N443_15 ( .fault(fault), .net(N443), .FEN(FEN[191]), .op(N443_t15) );
fim FAN_N460_0 ( .fault(fault), .net(N460), .FEN(FEN[192]), .op(N460_t0) );
fim FAN_N460_1 ( .fault(fault), .net(N460), .FEN(FEN[193]), .op(N460_t1) );
fim FAN_N460_2 ( .fault(fault), .net(N460), .FEN(FEN[194]), .op(N460_t2) );
fim FAN_N460_3 ( .fault(fault), .net(N460), .FEN(FEN[195]), .op(N460_t3) );
fim FAN_N460_4 ( .fault(fault), .net(N460), .FEN(FEN[196]), .op(N460_t4) );
fim FAN_N460_5 ( .fault(fault), .net(N460), .FEN(FEN[197]), .op(N460_t5) );
fim FAN_N460_6 ( .fault(fault), .net(N460), .FEN(FEN[198]), .op(N460_t6) );
fim FAN_N460_7 ( .fault(fault), .net(N460), .FEN(FEN[199]), .op(N460_t7) );
fim FAN_N460_8 ( .fault(fault), .net(N460), .FEN(FEN[200]), .op(N460_t8) );
fim FAN_N460_9 ( .fault(fault), .net(N460), .FEN(FEN[201]), .op(N460_t9) );
fim FAN_N460_10 ( .fault(fault), .net(N460), .FEN(FEN[202]), .op(N460_t10) );
fim FAN_N460_11 ( .fault(fault), .net(N460), .FEN(FEN[203]), .op(N460_t11) );
fim FAN_N460_12 ( .fault(fault), .net(N460), .FEN(FEN[204]), .op(N460_t12) );
fim FAN_N460_13 ( .fault(fault), .net(N460), .FEN(FEN[205]), .op(N460_t13) );
fim FAN_N460_14 ( .fault(fault), .net(N460), .FEN(FEN[206]), .op(N460_t14) );
fim FAN_N460_15 ( .fault(fault), .net(N460), .FEN(FEN[207]), .op(N460_t15) );
fim FAN_N477_0 ( .fault(fault), .net(N477), .FEN(FEN[208]), .op(N477_t0) );
fim FAN_N477_1 ( .fault(fault), .net(N477), .FEN(FEN[209]), .op(N477_t1) );
fim FAN_N477_2 ( .fault(fault), .net(N477), .FEN(FEN[210]), .op(N477_t2) );
fim FAN_N477_3 ( .fault(fault), .net(N477), .FEN(FEN[211]), .op(N477_t3) );
fim FAN_N477_4 ( .fault(fault), .net(N477), .FEN(FEN[212]), .op(N477_t4) );
fim FAN_N477_5 ( .fault(fault), .net(N477), .FEN(FEN[213]), .op(N477_t5) );
fim FAN_N477_6 ( .fault(fault), .net(N477), .FEN(FEN[214]), .op(N477_t6) );
fim FAN_N477_7 ( .fault(fault), .net(N477), .FEN(FEN[215]), .op(N477_t7) );
fim FAN_N477_8 ( .fault(fault), .net(N477), .FEN(FEN[216]), .op(N477_t8) );
fim FAN_N477_9 ( .fault(fault), .net(N477), .FEN(FEN[217]), .op(N477_t9) );
fim FAN_N477_10 ( .fault(fault), .net(N477), .FEN(FEN[218]), .op(N477_t10) );
fim FAN_N477_11 ( .fault(fault), .net(N477), .FEN(FEN[219]), .op(N477_t11) );
fim FAN_N477_12 ( .fault(fault), .net(N477), .FEN(FEN[220]), .op(N477_t12) );
fim FAN_N477_13 ( .fault(fault), .net(N477), .FEN(FEN[221]), .op(N477_t13) );
fim FAN_N477_14 ( .fault(fault), .net(N477), .FEN(FEN[222]), .op(N477_t14) );
fim FAN_N477_15 ( .fault(fault), .net(N477), .FEN(FEN[223]), .op(N477_t15) );
fim FAN_N494_0 ( .fault(fault), .net(N494), .FEN(FEN[224]), .op(N494_t0) );
fim FAN_N494_1 ( .fault(fault), .net(N494), .FEN(FEN[225]), .op(N494_t1) );
fim FAN_N494_2 ( .fault(fault), .net(N494), .FEN(FEN[226]), .op(N494_t2) );
fim FAN_N494_3 ( .fault(fault), .net(N494), .FEN(FEN[227]), .op(N494_t3) );
fim FAN_N494_4 ( .fault(fault), .net(N494), .FEN(FEN[228]), .op(N494_t4) );
fim FAN_N494_5 ( .fault(fault), .net(N494), .FEN(FEN[229]), .op(N494_t5) );
fim FAN_N494_6 ( .fault(fault), .net(N494), .FEN(FEN[230]), .op(N494_t6) );
fim FAN_N494_7 ( .fault(fault), .net(N494), .FEN(FEN[231]), .op(N494_t7) );
fim FAN_N494_8 ( .fault(fault), .net(N494), .FEN(FEN[232]), .op(N494_t8) );
fim FAN_N494_9 ( .fault(fault), .net(N494), .FEN(FEN[233]), .op(N494_t9) );
fim FAN_N494_10 ( .fault(fault), .net(N494), .FEN(FEN[234]), .op(N494_t10) );
fim FAN_N494_11 ( .fault(fault), .net(N494), .FEN(FEN[235]), .op(N494_t11) );
fim FAN_N494_12 ( .fault(fault), .net(N494), .FEN(FEN[236]), .op(N494_t12) );
fim FAN_N494_13 ( .fault(fault), .net(N494), .FEN(FEN[237]), .op(N494_t13) );
fim FAN_N494_14 ( .fault(fault), .net(N494), .FEN(FEN[238]), .op(N494_t14) );
fim FAN_N494_15 ( .fault(fault), .net(N494), .FEN(FEN[239]), .op(N494_t15) );
fim FAN_N511_0 ( .fault(fault), .net(N511), .FEN(FEN[240]), .op(N511_t0) );
fim FAN_N511_1 ( .fault(fault), .net(N511), .FEN(FEN[241]), .op(N511_t1) );
fim FAN_N511_2 ( .fault(fault), .net(N511), .FEN(FEN[242]), .op(N511_t2) );
fim FAN_N511_3 ( .fault(fault), .net(N511), .FEN(FEN[243]), .op(N511_t3) );
fim FAN_N511_4 ( .fault(fault), .net(N511), .FEN(FEN[244]), .op(N511_t4) );
fim FAN_N511_5 ( .fault(fault), .net(N511), .FEN(FEN[245]), .op(N511_t5) );
fim FAN_N511_6 ( .fault(fault), .net(N511), .FEN(FEN[246]), .op(N511_t6) );
fim FAN_N511_7 ( .fault(fault), .net(N511), .FEN(FEN[247]), .op(N511_t7) );
fim FAN_N511_8 ( .fault(fault), .net(N511), .FEN(FEN[248]), .op(N511_t8) );
fim FAN_N511_9 ( .fault(fault), .net(N511), .FEN(FEN[249]), .op(N511_t9) );
fim FAN_N511_10 ( .fault(fault), .net(N511), .FEN(FEN[250]), .op(N511_t10) );
fim FAN_N511_11 ( .fault(fault), .net(N511), .FEN(FEN[251]), .op(N511_t11) );
fim FAN_N511_12 ( .fault(fault), .net(N511), .FEN(FEN[252]), .op(N511_t12) );
fim FAN_N511_13 ( .fault(fault), .net(N511), .FEN(FEN[253]), .op(N511_t13) );
fim FAN_N511_14 ( .fault(fault), .net(N511), .FEN(FEN[254]), .op(N511_t14) );
fim FAN_N511_15 ( .fault(fault), .net(N511), .FEN(FEN[255]), .op(N511_t15) );
fim FAN_N528_0 ( .fault(fault), .net(N528), .FEN(FEN[256]), .op(N528_t0) );
fim FAN_N528_1 ( .fault(fault), .net(N528), .FEN(FEN[257]), .op(N528_t1) );
fim FAN_N528_2 ( .fault(fault), .net(N528), .FEN(FEN[258]), .op(N528_t2) );
fim FAN_N528_3 ( .fault(fault), .net(N528), .FEN(FEN[259]), .op(N528_t3) );
fim FAN_N528_4 ( .fault(fault), .net(N528), .FEN(FEN[260]), .op(N528_t4) );
fim FAN_N528_5 ( .fault(fault), .net(N528), .FEN(FEN[261]), .op(N528_t5) );
fim FAN_N528_6 ( .fault(fault), .net(N528), .FEN(FEN[262]), .op(N528_t6) );
fim FAN_N528_7 ( .fault(fault), .net(N528), .FEN(FEN[263]), .op(N528_t7) );
fim FAN_N528_8 ( .fault(fault), .net(N528), .FEN(FEN[264]), .op(N528_t8) );
fim FAN_N528_9 ( .fault(fault), .net(N528), .FEN(FEN[265]), .op(N528_t9) );
fim FAN_N528_10 ( .fault(fault), .net(N528), .FEN(FEN[266]), .op(N528_t10) );
fim FAN_N528_11 ( .fault(fault), .net(N528), .FEN(FEN[267]), .op(N528_t11) );
fim FAN_N528_12 ( .fault(fault), .net(N528), .FEN(FEN[268]), .op(N528_t12) );
fim FAN_N528_13 ( .fault(fault), .net(N528), .FEN(FEN[269]), .op(N528_t13) );
fim FAN_N528_14 ( .fault(fault), .net(N528), .FEN(FEN[270]), .op(N528_t14) );
fim FAN_N528_15 ( .fault(fault), .net(N528), .FEN(FEN[271]), .op(N528_t15) );
fim FAN_N18_0 ( .fault(fault), .net(N18), .FEN(FEN[272]), .op(N18_t0) );
fim FAN_N18_1 ( .fault(fault), .net(N18), .FEN(FEN[273]), .op(N18_t1) );
fim FAN_N18_2 ( .fault(fault), .net(N18), .FEN(FEN[274]), .op(N18_t2) );
fim FAN_N18_3 ( .fault(fault), .net(N18), .FEN(FEN[275]), .op(N18_t3) );
fim FAN_N18_4 ( .fault(fault), .net(N18), .FEN(FEN[276]), .op(N18_t4) );
fim FAN_N18_5 ( .fault(fault), .net(N18), .FEN(FEN[277]), .op(N18_t5) );
fim FAN_N18_6 ( .fault(fault), .net(N18), .FEN(FEN[278]), .op(N18_t6) );
fim FAN_N18_7 ( .fault(fault), .net(N18), .FEN(FEN[279]), .op(N18_t7) );
fim FAN_N18_8 ( .fault(fault), .net(N18), .FEN(FEN[280]), .op(N18_t8) );
fim FAN_N18_9 ( .fault(fault), .net(N18), .FEN(FEN[281]), .op(N18_t9) );
fim FAN_N18_10 ( .fault(fault), .net(N18), .FEN(FEN[282]), .op(N18_t10) );
fim FAN_N18_11 ( .fault(fault), .net(N18), .FEN(FEN[283]), .op(N18_t11) );
fim FAN_N18_12 ( .fault(fault), .net(N18), .FEN(FEN[284]), .op(N18_t12) );
fim FAN_N18_13 ( .fault(fault), .net(N18), .FEN(FEN[285]), .op(N18_t13) );
fim FAN_N18_14 ( .fault(fault), .net(N18), .FEN(FEN[286]), .op(N18_t14) );
fim FAN_N18_15 ( .fault(fault), .net(N18), .FEN(FEN[287]), .op(N18_t15) );
fim FAN_N35_0 ( .fault(fault), .net(N35), .FEN(FEN[288]), .op(N35_t0) );
fim FAN_N35_1 ( .fault(fault), .net(N35), .FEN(FEN[289]), .op(N35_t1) );
fim FAN_N35_2 ( .fault(fault), .net(N35), .FEN(FEN[290]), .op(N35_t2) );
fim FAN_N35_3 ( .fault(fault), .net(N35), .FEN(FEN[291]), .op(N35_t3) );
fim FAN_N35_4 ( .fault(fault), .net(N35), .FEN(FEN[292]), .op(N35_t4) );
fim FAN_N35_5 ( .fault(fault), .net(N35), .FEN(FEN[293]), .op(N35_t5) );
fim FAN_N35_6 ( .fault(fault), .net(N35), .FEN(FEN[294]), .op(N35_t6) );
fim FAN_N35_7 ( .fault(fault), .net(N35), .FEN(FEN[295]), .op(N35_t7) );
fim FAN_N35_8 ( .fault(fault), .net(N35), .FEN(FEN[296]), .op(N35_t8) );
fim FAN_N35_9 ( .fault(fault), .net(N35), .FEN(FEN[297]), .op(N35_t9) );
fim FAN_N35_10 ( .fault(fault), .net(N35), .FEN(FEN[298]), .op(N35_t10) );
fim FAN_N35_11 ( .fault(fault), .net(N35), .FEN(FEN[299]), .op(N35_t11) );
fim FAN_N35_12 ( .fault(fault), .net(N35), .FEN(FEN[300]), .op(N35_t12) );
fim FAN_N35_13 ( .fault(fault), .net(N35), .FEN(FEN[301]), .op(N35_t13) );
fim FAN_N35_14 ( .fault(fault), .net(N35), .FEN(FEN[302]), .op(N35_t14) );
fim FAN_N35_15 ( .fault(fault), .net(N35), .FEN(FEN[303]), .op(N35_t15) );
fim FAN_N52_0 ( .fault(fault), .net(N52), .FEN(FEN[304]), .op(N52_t0) );
fim FAN_N52_1 ( .fault(fault), .net(N52), .FEN(FEN[305]), .op(N52_t1) );
fim FAN_N52_2 ( .fault(fault), .net(N52), .FEN(FEN[306]), .op(N52_t2) );
fim FAN_N52_3 ( .fault(fault), .net(N52), .FEN(FEN[307]), .op(N52_t3) );
fim FAN_N52_4 ( .fault(fault), .net(N52), .FEN(FEN[308]), .op(N52_t4) );
fim FAN_N52_5 ( .fault(fault), .net(N52), .FEN(FEN[309]), .op(N52_t5) );
fim FAN_N52_6 ( .fault(fault), .net(N52), .FEN(FEN[310]), .op(N52_t6) );
fim FAN_N52_7 ( .fault(fault), .net(N52), .FEN(FEN[311]), .op(N52_t7) );
fim FAN_N52_8 ( .fault(fault), .net(N52), .FEN(FEN[312]), .op(N52_t8) );
fim FAN_N52_9 ( .fault(fault), .net(N52), .FEN(FEN[313]), .op(N52_t9) );
fim FAN_N52_10 ( .fault(fault), .net(N52), .FEN(FEN[314]), .op(N52_t10) );
fim FAN_N52_11 ( .fault(fault), .net(N52), .FEN(FEN[315]), .op(N52_t11) );
fim FAN_N52_12 ( .fault(fault), .net(N52), .FEN(FEN[316]), .op(N52_t12) );
fim FAN_N52_13 ( .fault(fault), .net(N52), .FEN(FEN[317]), .op(N52_t13) );
fim FAN_N52_14 ( .fault(fault), .net(N52), .FEN(FEN[318]), .op(N52_t14) );
fim FAN_N52_15 ( .fault(fault), .net(N52), .FEN(FEN[319]), .op(N52_t15) );
fim FAN_N69_0 ( .fault(fault), .net(N69), .FEN(FEN[320]), .op(N69_t0) );
fim FAN_N69_1 ( .fault(fault), .net(N69), .FEN(FEN[321]), .op(N69_t1) );
fim FAN_N69_2 ( .fault(fault), .net(N69), .FEN(FEN[322]), .op(N69_t2) );
fim FAN_N69_3 ( .fault(fault), .net(N69), .FEN(FEN[323]), .op(N69_t3) );
fim FAN_N69_4 ( .fault(fault), .net(N69), .FEN(FEN[324]), .op(N69_t4) );
fim FAN_N69_5 ( .fault(fault), .net(N69), .FEN(FEN[325]), .op(N69_t5) );
fim FAN_N69_6 ( .fault(fault), .net(N69), .FEN(FEN[326]), .op(N69_t6) );
fim FAN_N69_7 ( .fault(fault), .net(N69), .FEN(FEN[327]), .op(N69_t7) );
fim FAN_N69_8 ( .fault(fault), .net(N69), .FEN(FEN[328]), .op(N69_t8) );
fim FAN_N69_9 ( .fault(fault), .net(N69), .FEN(FEN[329]), .op(N69_t9) );
fim FAN_N69_10 ( .fault(fault), .net(N69), .FEN(FEN[330]), .op(N69_t10) );
fim FAN_N69_11 ( .fault(fault), .net(N69), .FEN(FEN[331]), .op(N69_t11) );
fim FAN_N69_12 ( .fault(fault), .net(N69), .FEN(FEN[332]), .op(N69_t12) );
fim FAN_N69_13 ( .fault(fault), .net(N69), .FEN(FEN[333]), .op(N69_t13) );
fim FAN_N69_14 ( .fault(fault), .net(N69), .FEN(FEN[334]), .op(N69_t14) );
fim FAN_N69_15 ( .fault(fault), .net(N69), .FEN(FEN[335]), .op(N69_t15) );
fim FAN_N86_0 ( .fault(fault), .net(N86), .FEN(FEN[336]), .op(N86_t0) );
fim FAN_N86_1 ( .fault(fault), .net(N86), .FEN(FEN[337]), .op(N86_t1) );
fim FAN_N86_2 ( .fault(fault), .net(N86), .FEN(FEN[338]), .op(N86_t2) );
fim FAN_N86_3 ( .fault(fault), .net(N86), .FEN(FEN[339]), .op(N86_t3) );
fim FAN_N86_4 ( .fault(fault), .net(N86), .FEN(FEN[340]), .op(N86_t4) );
fim FAN_N86_5 ( .fault(fault), .net(N86), .FEN(FEN[341]), .op(N86_t5) );
fim FAN_N86_6 ( .fault(fault), .net(N86), .FEN(FEN[342]), .op(N86_t6) );
fim FAN_N86_7 ( .fault(fault), .net(N86), .FEN(FEN[343]), .op(N86_t7) );
fim FAN_N86_8 ( .fault(fault), .net(N86), .FEN(FEN[344]), .op(N86_t8) );
fim FAN_N86_9 ( .fault(fault), .net(N86), .FEN(FEN[345]), .op(N86_t9) );
fim FAN_N86_10 ( .fault(fault), .net(N86), .FEN(FEN[346]), .op(N86_t10) );
fim FAN_N86_11 ( .fault(fault), .net(N86), .FEN(FEN[347]), .op(N86_t11) );
fim FAN_N86_12 ( .fault(fault), .net(N86), .FEN(FEN[348]), .op(N86_t12) );
fim FAN_N86_13 ( .fault(fault), .net(N86), .FEN(FEN[349]), .op(N86_t13) );
fim FAN_N86_14 ( .fault(fault), .net(N86), .FEN(FEN[350]), .op(N86_t14) );
fim FAN_N86_15 ( .fault(fault), .net(N86), .FEN(FEN[351]), .op(N86_t15) );
fim FAN_N103_0 ( .fault(fault), .net(N103), .FEN(FEN[352]), .op(N103_t0) );
fim FAN_N103_1 ( .fault(fault), .net(N103), .FEN(FEN[353]), .op(N103_t1) );
fim FAN_N103_2 ( .fault(fault), .net(N103), .FEN(FEN[354]), .op(N103_t2) );
fim FAN_N103_3 ( .fault(fault), .net(N103), .FEN(FEN[355]), .op(N103_t3) );
fim FAN_N103_4 ( .fault(fault), .net(N103), .FEN(FEN[356]), .op(N103_t4) );
fim FAN_N103_5 ( .fault(fault), .net(N103), .FEN(FEN[357]), .op(N103_t5) );
fim FAN_N103_6 ( .fault(fault), .net(N103), .FEN(FEN[358]), .op(N103_t6) );
fim FAN_N103_7 ( .fault(fault), .net(N103), .FEN(FEN[359]), .op(N103_t7) );
fim FAN_N103_8 ( .fault(fault), .net(N103), .FEN(FEN[360]), .op(N103_t8) );
fim FAN_N103_9 ( .fault(fault), .net(N103), .FEN(FEN[361]), .op(N103_t9) );
fim FAN_N103_10 ( .fault(fault), .net(N103), .FEN(FEN[362]), .op(N103_t10) );
fim FAN_N103_11 ( .fault(fault), .net(N103), .FEN(FEN[363]), .op(N103_t11) );
fim FAN_N103_12 ( .fault(fault), .net(N103), .FEN(FEN[364]), .op(N103_t12) );
fim FAN_N103_13 ( .fault(fault), .net(N103), .FEN(FEN[365]), .op(N103_t13) );
fim FAN_N103_14 ( .fault(fault), .net(N103), .FEN(FEN[366]), .op(N103_t14) );
fim FAN_N103_15 ( .fault(fault), .net(N103), .FEN(FEN[367]), .op(N103_t15) );
fim FAN_N120_0 ( .fault(fault), .net(N120), .FEN(FEN[368]), .op(N120_t0) );
fim FAN_N120_1 ( .fault(fault), .net(N120), .FEN(FEN[369]), .op(N120_t1) );
fim FAN_N120_2 ( .fault(fault), .net(N120), .FEN(FEN[370]), .op(N120_t2) );
fim FAN_N120_3 ( .fault(fault), .net(N120), .FEN(FEN[371]), .op(N120_t3) );
fim FAN_N120_4 ( .fault(fault), .net(N120), .FEN(FEN[372]), .op(N120_t4) );
fim FAN_N120_5 ( .fault(fault), .net(N120), .FEN(FEN[373]), .op(N120_t5) );
fim FAN_N120_6 ( .fault(fault), .net(N120), .FEN(FEN[374]), .op(N120_t6) );
fim FAN_N120_7 ( .fault(fault), .net(N120), .FEN(FEN[375]), .op(N120_t7) );
fim FAN_N120_8 ( .fault(fault), .net(N120), .FEN(FEN[376]), .op(N120_t8) );
fim FAN_N120_9 ( .fault(fault), .net(N120), .FEN(FEN[377]), .op(N120_t9) );
fim FAN_N120_10 ( .fault(fault), .net(N120), .FEN(FEN[378]), .op(N120_t10) );
fim FAN_N120_11 ( .fault(fault), .net(N120), .FEN(FEN[379]), .op(N120_t11) );
fim FAN_N120_12 ( .fault(fault), .net(N120), .FEN(FEN[380]), .op(N120_t12) );
fim FAN_N120_13 ( .fault(fault), .net(N120), .FEN(FEN[381]), .op(N120_t13) );
fim FAN_N120_14 ( .fault(fault), .net(N120), .FEN(FEN[382]), .op(N120_t14) );
fim FAN_N120_15 ( .fault(fault), .net(N120), .FEN(FEN[383]), .op(N120_t15) );
fim FAN_N137_0 ( .fault(fault), .net(N137), .FEN(FEN[384]), .op(N137_t0) );
fim FAN_N137_1 ( .fault(fault), .net(N137), .FEN(FEN[385]), .op(N137_t1) );
fim FAN_N137_2 ( .fault(fault), .net(N137), .FEN(FEN[386]), .op(N137_t2) );
fim FAN_N137_3 ( .fault(fault), .net(N137), .FEN(FEN[387]), .op(N137_t3) );
fim FAN_N137_4 ( .fault(fault), .net(N137), .FEN(FEN[388]), .op(N137_t4) );
fim FAN_N137_5 ( .fault(fault), .net(N137), .FEN(FEN[389]), .op(N137_t5) );
fim FAN_N137_6 ( .fault(fault), .net(N137), .FEN(FEN[390]), .op(N137_t6) );
fim FAN_N137_7 ( .fault(fault), .net(N137), .FEN(FEN[391]), .op(N137_t7) );
fim FAN_N137_8 ( .fault(fault), .net(N137), .FEN(FEN[392]), .op(N137_t8) );
fim FAN_N137_9 ( .fault(fault), .net(N137), .FEN(FEN[393]), .op(N137_t9) );
fim FAN_N137_10 ( .fault(fault), .net(N137), .FEN(FEN[394]), .op(N137_t10) );
fim FAN_N137_11 ( .fault(fault), .net(N137), .FEN(FEN[395]), .op(N137_t11) );
fim FAN_N137_12 ( .fault(fault), .net(N137), .FEN(FEN[396]), .op(N137_t12) );
fim FAN_N137_13 ( .fault(fault), .net(N137), .FEN(FEN[397]), .op(N137_t13) );
fim FAN_N137_14 ( .fault(fault), .net(N137), .FEN(FEN[398]), .op(N137_t14) );
fim FAN_N137_15 ( .fault(fault), .net(N137), .FEN(FEN[399]), .op(N137_t15) );
fim FAN_N154_0 ( .fault(fault), .net(N154), .FEN(FEN[400]), .op(N154_t0) );
fim FAN_N154_1 ( .fault(fault), .net(N154), .FEN(FEN[401]), .op(N154_t1) );
fim FAN_N154_2 ( .fault(fault), .net(N154), .FEN(FEN[402]), .op(N154_t2) );
fim FAN_N154_3 ( .fault(fault), .net(N154), .FEN(FEN[403]), .op(N154_t3) );
fim FAN_N154_4 ( .fault(fault), .net(N154), .FEN(FEN[404]), .op(N154_t4) );
fim FAN_N154_5 ( .fault(fault), .net(N154), .FEN(FEN[405]), .op(N154_t5) );
fim FAN_N154_6 ( .fault(fault), .net(N154), .FEN(FEN[406]), .op(N154_t6) );
fim FAN_N154_7 ( .fault(fault), .net(N154), .FEN(FEN[407]), .op(N154_t7) );
fim FAN_N154_8 ( .fault(fault), .net(N154), .FEN(FEN[408]), .op(N154_t8) );
fim FAN_N154_9 ( .fault(fault), .net(N154), .FEN(FEN[409]), .op(N154_t9) );
fim FAN_N154_10 ( .fault(fault), .net(N154), .FEN(FEN[410]), .op(N154_t10) );
fim FAN_N154_11 ( .fault(fault), .net(N154), .FEN(FEN[411]), .op(N154_t11) );
fim FAN_N154_12 ( .fault(fault), .net(N154), .FEN(FEN[412]), .op(N154_t12) );
fim FAN_N154_13 ( .fault(fault), .net(N154), .FEN(FEN[413]), .op(N154_t13) );
fim FAN_N154_14 ( .fault(fault), .net(N154), .FEN(FEN[414]), .op(N154_t14) );
fim FAN_N154_15 ( .fault(fault), .net(N154), .FEN(FEN[415]), .op(N154_t15) );
fim FAN_N171_0 ( .fault(fault), .net(N171), .FEN(FEN[416]), .op(N171_t0) );
fim FAN_N171_1 ( .fault(fault), .net(N171), .FEN(FEN[417]), .op(N171_t1) );
fim FAN_N171_2 ( .fault(fault), .net(N171), .FEN(FEN[418]), .op(N171_t2) );
fim FAN_N171_3 ( .fault(fault), .net(N171), .FEN(FEN[419]), .op(N171_t3) );
fim FAN_N171_4 ( .fault(fault), .net(N171), .FEN(FEN[420]), .op(N171_t4) );
fim FAN_N171_5 ( .fault(fault), .net(N171), .FEN(FEN[421]), .op(N171_t5) );
fim FAN_N171_6 ( .fault(fault), .net(N171), .FEN(FEN[422]), .op(N171_t6) );
fim FAN_N171_7 ( .fault(fault), .net(N171), .FEN(FEN[423]), .op(N171_t7) );
fim FAN_N171_8 ( .fault(fault), .net(N171), .FEN(FEN[424]), .op(N171_t8) );
fim FAN_N171_9 ( .fault(fault), .net(N171), .FEN(FEN[425]), .op(N171_t9) );
fim FAN_N171_10 ( .fault(fault), .net(N171), .FEN(FEN[426]), .op(N171_t10) );
fim FAN_N171_11 ( .fault(fault), .net(N171), .FEN(FEN[427]), .op(N171_t11) );
fim FAN_N171_12 ( .fault(fault), .net(N171), .FEN(FEN[428]), .op(N171_t12) );
fim FAN_N171_13 ( .fault(fault), .net(N171), .FEN(FEN[429]), .op(N171_t13) );
fim FAN_N171_14 ( .fault(fault), .net(N171), .FEN(FEN[430]), .op(N171_t14) );
fim FAN_N171_15 ( .fault(fault), .net(N171), .FEN(FEN[431]), .op(N171_t15) );
fim FAN_N188_0 ( .fault(fault), .net(N188), .FEN(FEN[432]), .op(N188_t0) );
fim FAN_N188_1 ( .fault(fault), .net(N188), .FEN(FEN[433]), .op(N188_t1) );
fim FAN_N188_2 ( .fault(fault), .net(N188), .FEN(FEN[434]), .op(N188_t2) );
fim FAN_N188_3 ( .fault(fault), .net(N188), .FEN(FEN[435]), .op(N188_t3) );
fim FAN_N188_4 ( .fault(fault), .net(N188), .FEN(FEN[436]), .op(N188_t4) );
fim FAN_N188_5 ( .fault(fault), .net(N188), .FEN(FEN[437]), .op(N188_t5) );
fim FAN_N188_6 ( .fault(fault), .net(N188), .FEN(FEN[438]), .op(N188_t6) );
fim FAN_N188_7 ( .fault(fault), .net(N188), .FEN(FEN[439]), .op(N188_t7) );
fim FAN_N188_8 ( .fault(fault), .net(N188), .FEN(FEN[440]), .op(N188_t8) );
fim FAN_N188_9 ( .fault(fault), .net(N188), .FEN(FEN[441]), .op(N188_t9) );
fim FAN_N188_10 ( .fault(fault), .net(N188), .FEN(FEN[442]), .op(N188_t10) );
fim FAN_N188_11 ( .fault(fault), .net(N188), .FEN(FEN[443]), .op(N188_t11) );
fim FAN_N188_12 ( .fault(fault), .net(N188), .FEN(FEN[444]), .op(N188_t12) );
fim FAN_N188_13 ( .fault(fault), .net(N188), .FEN(FEN[445]), .op(N188_t13) );
fim FAN_N188_14 ( .fault(fault), .net(N188), .FEN(FEN[446]), .op(N188_t14) );
fim FAN_N188_15 ( .fault(fault), .net(N188), .FEN(FEN[447]), .op(N188_t15) );
fim FAN_N205_0 ( .fault(fault), .net(N205), .FEN(FEN[448]), .op(N205_t0) );
fim FAN_N205_1 ( .fault(fault), .net(N205), .FEN(FEN[449]), .op(N205_t1) );
fim FAN_N205_2 ( .fault(fault), .net(N205), .FEN(FEN[450]), .op(N205_t2) );
fim FAN_N205_3 ( .fault(fault), .net(N205), .FEN(FEN[451]), .op(N205_t3) );
fim FAN_N205_4 ( .fault(fault), .net(N205), .FEN(FEN[452]), .op(N205_t4) );
fim FAN_N205_5 ( .fault(fault), .net(N205), .FEN(FEN[453]), .op(N205_t5) );
fim FAN_N205_6 ( .fault(fault), .net(N205), .FEN(FEN[454]), .op(N205_t6) );
fim FAN_N205_7 ( .fault(fault), .net(N205), .FEN(FEN[455]), .op(N205_t7) );
fim FAN_N205_8 ( .fault(fault), .net(N205), .FEN(FEN[456]), .op(N205_t8) );
fim FAN_N205_9 ( .fault(fault), .net(N205), .FEN(FEN[457]), .op(N205_t9) );
fim FAN_N205_10 ( .fault(fault), .net(N205), .FEN(FEN[458]), .op(N205_t10) );
fim FAN_N205_11 ( .fault(fault), .net(N205), .FEN(FEN[459]), .op(N205_t11) );
fim FAN_N205_12 ( .fault(fault), .net(N205), .FEN(FEN[460]), .op(N205_t12) );
fim FAN_N205_13 ( .fault(fault), .net(N205), .FEN(FEN[461]), .op(N205_t13) );
fim FAN_N205_14 ( .fault(fault), .net(N205), .FEN(FEN[462]), .op(N205_t14) );
fim FAN_N205_15 ( .fault(fault), .net(N205), .FEN(FEN[463]), .op(N205_t15) );
fim FAN_N222_0 ( .fault(fault), .net(N222), .FEN(FEN[464]), .op(N222_t0) );
fim FAN_N222_1 ( .fault(fault), .net(N222), .FEN(FEN[465]), .op(N222_t1) );
fim FAN_N222_2 ( .fault(fault), .net(N222), .FEN(FEN[466]), .op(N222_t2) );
fim FAN_N222_3 ( .fault(fault), .net(N222), .FEN(FEN[467]), .op(N222_t3) );
fim FAN_N222_4 ( .fault(fault), .net(N222), .FEN(FEN[468]), .op(N222_t4) );
fim FAN_N222_5 ( .fault(fault), .net(N222), .FEN(FEN[469]), .op(N222_t5) );
fim FAN_N222_6 ( .fault(fault), .net(N222), .FEN(FEN[470]), .op(N222_t6) );
fim FAN_N222_7 ( .fault(fault), .net(N222), .FEN(FEN[471]), .op(N222_t7) );
fim FAN_N222_8 ( .fault(fault), .net(N222), .FEN(FEN[472]), .op(N222_t8) );
fim FAN_N222_9 ( .fault(fault), .net(N222), .FEN(FEN[473]), .op(N222_t9) );
fim FAN_N222_10 ( .fault(fault), .net(N222), .FEN(FEN[474]), .op(N222_t10) );
fim FAN_N222_11 ( .fault(fault), .net(N222), .FEN(FEN[475]), .op(N222_t11) );
fim FAN_N222_12 ( .fault(fault), .net(N222), .FEN(FEN[476]), .op(N222_t12) );
fim FAN_N222_13 ( .fault(fault), .net(N222), .FEN(FEN[477]), .op(N222_t13) );
fim FAN_N222_14 ( .fault(fault), .net(N222), .FEN(FEN[478]), .op(N222_t14) );
fim FAN_N222_15 ( .fault(fault), .net(N222), .FEN(FEN[479]), .op(N222_t15) );
fim FAN_N239_0 ( .fault(fault), .net(N239), .FEN(FEN[480]), .op(N239_t0) );
fim FAN_N239_1 ( .fault(fault), .net(N239), .FEN(FEN[481]), .op(N239_t1) );
fim FAN_N239_2 ( .fault(fault), .net(N239), .FEN(FEN[482]), .op(N239_t2) );
fim FAN_N239_3 ( .fault(fault), .net(N239), .FEN(FEN[483]), .op(N239_t3) );
fim FAN_N239_4 ( .fault(fault), .net(N239), .FEN(FEN[484]), .op(N239_t4) );
fim FAN_N239_5 ( .fault(fault), .net(N239), .FEN(FEN[485]), .op(N239_t5) );
fim FAN_N239_6 ( .fault(fault), .net(N239), .FEN(FEN[486]), .op(N239_t6) );
fim FAN_N239_7 ( .fault(fault), .net(N239), .FEN(FEN[487]), .op(N239_t7) );
fim FAN_N239_8 ( .fault(fault), .net(N239), .FEN(FEN[488]), .op(N239_t8) );
fim FAN_N239_9 ( .fault(fault), .net(N239), .FEN(FEN[489]), .op(N239_t9) );
fim FAN_N239_10 ( .fault(fault), .net(N239), .FEN(FEN[490]), .op(N239_t10) );
fim FAN_N239_11 ( .fault(fault), .net(N239), .FEN(FEN[491]), .op(N239_t11) );
fim FAN_N239_12 ( .fault(fault), .net(N239), .FEN(FEN[492]), .op(N239_t12) );
fim FAN_N239_13 ( .fault(fault), .net(N239), .FEN(FEN[493]), .op(N239_t13) );
fim FAN_N239_14 ( .fault(fault), .net(N239), .FEN(FEN[494]), .op(N239_t14) );
fim FAN_N239_15 ( .fault(fault), .net(N239), .FEN(FEN[495]), .op(N239_t15) );
fim FAN_N256_0 ( .fault(fault), .net(N256), .FEN(FEN[496]), .op(N256_t0) );
fim FAN_N256_1 ( .fault(fault), .net(N256), .FEN(FEN[497]), .op(N256_t1) );
fim FAN_N256_2 ( .fault(fault), .net(N256), .FEN(FEN[498]), .op(N256_t2) );
fim FAN_N256_3 ( .fault(fault), .net(N256), .FEN(FEN[499]), .op(N256_t3) );
fim FAN_N256_4 ( .fault(fault), .net(N256), .FEN(FEN[500]), .op(N256_t4) );
fim FAN_N256_5 ( .fault(fault), .net(N256), .FEN(FEN[501]), .op(N256_t5) );
fim FAN_N256_6 ( .fault(fault), .net(N256), .FEN(FEN[502]), .op(N256_t6) );
fim FAN_N256_7 ( .fault(fault), .net(N256), .FEN(FEN[503]), .op(N256_t7) );
fim FAN_N256_8 ( .fault(fault), .net(N256), .FEN(FEN[504]), .op(N256_t8) );
fim FAN_N256_9 ( .fault(fault), .net(N256), .FEN(FEN[505]), .op(N256_t9) );
fim FAN_N256_10 ( .fault(fault), .net(N256), .FEN(FEN[506]), .op(N256_t10) );
fim FAN_N256_11 ( .fault(fault), .net(N256), .FEN(FEN[507]), .op(N256_t11) );
fim FAN_N256_12 ( .fault(fault), .net(N256), .FEN(FEN[508]), .op(N256_t12) );
fim FAN_N256_13 ( .fault(fault), .net(N256), .FEN(FEN[509]), .op(N256_t13) );
fim FAN_N256_14 ( .fault(fault), .net(N256), .FEN(FEN[510]), .op(N256_t14) );
fim FAN_N256_15 ( .fault(fault), .net(N256), .FEN(FEN[511]), .op(N256_t15) );
fim FAN_N591_0 ( .fault(fault), .net(N591), .FEN(FEN[512]), .op(N591_t0) );
fim FAN_N591_1 ( .fault(fault), .net(N591), .FEN(FEN[513]), .op(N591_t1) );
fim FAN_N639_0 ( .fault(fault), .net(N639), .FEN(FEN[514]), .op(N639_t0) );
fim FAN_N639_1 ( .fault(fault), .net(N639), .FEN(FEN[515]), .op(N639_t1) );
fim FAN_N687_0 ( .fault(fault), .net(N687), .FEN(FEN[516]), .op(N687_t0) );
fim FAN_N687_1 ( .fault(fault), .net(N687), .FEN(FEN[517]), .op(N687_t1) );
fim FAN_N735_0 ( .fault(fault), .net(N735), .FEN(FEN[518]), .op(N735_t0) );
fim FAN_N735_1 ( .fault(fault), .net(N735), .FEN(FEN[519]), .op(N735_t1) );
fim FAN_N783_0 ( .fault(fault), .net(N783), .FEN(FEN[520]), .op(N783_t0) );
fim FAN_N783_1 ( .fault(fault), .net(N783), .FEN(FEN[521]), .op(N783_t1) );
fim FAN_N831_0 ( .fault(fault), .net(N831), .FEN(FEN[522]), .op(N831_t0) );
fim FAN_N831_1 ( .fault(fault), .net(N831), .FEN(FEN[523]), .op(N831_t1) );
fim FAN_N879_0 ( .fault(fault), .net(N879), .FEN(FEN[524]), .op(N879_t0) );
fim FAN_N879_1 ( .fault(fault), .net(N879), .FEN(FEN[525]), .op(N879_t1) );
fim FAN_N927_0 ( .fault(fault), .net(N927), .FEN(FEN[526]), .op(N927_t0) );
fim FAN_N927_1 ( .fault(fault), .net(N927), .FEN(FEN[527]), .op(N927_t1) );
fim FAN_N975_0 ( .fault(fault), .net(N975), .FEN(FEN[528]), .op(N975_t0) );
fim FAN_N975_1 ( .fault(fault), .net(N975), .FEN(FEN[529]), .op(N975_t1) );
fim FAN_N1023_0 ( .fault(fault), .net(N1023), .FEN(FEN[530]), .op(N1023_t0) );
fim FAN_N1023_1 ( .fault(fault), .net(N1023), .FEN(FEN[531]), .op(N1023_t1) );
fim FAN_N1071_0 ( .fault(fault), .net(N1071), .FEN(FEN[532]), .op(N1071_t0) );
fim FAN_N1071_1 ( .fault(fault), .net(N1071), .FEN(FEN[533]), .op(N1071_t1) );
fim FAN_N1119_0 ( .fault(fault), .net(N1119), .FEN(FEN[534]), .op(N1119_t0) );
fim FAN_N1119_1 ( .fault(fault), .net(N1119), .FEN(FEN[535]), .op(N1119_t1) );
fim FAN_N1167_0 ( .fault(fault), .net(N1167), .FEN(FEN[536]), .op(N1167_t0) );
fim FAN_N1167_1 ( .fault(fault), .net(N1167), .FEN(FEN[537]), .op(N1167_t1) );
fim FAN_N1215_0 ( .fault(fault), .net(N1215), .FEN(FEN[538]), .op(N1215_t0) );
fim FAN_N1215_1 ( .fault(fault), .net(N1215), .FEN(FEN[539]), .op(N1215_t1) );
fim FAN_N1263_0 ( .fault(fault), .net(N1263), .FEN(FEN[540]), .op(N1263_t0) );
fim FAN_N1263_1 ( .fault(fault), .net(N1263), .FEN(FEN[541]), .op(N1263_t1) );
fim FAN_N1311_0 ( .fault(fault), .net(N1311), .FEN(FEN[542]), .op(N1311_t0) );
fim FAN_N1311_1 ( .fault(fault), .net(N1311), .FEN(FEN[543]), .op(N1311_t1) );
fim FAN_N1311_2 ( .fault(fault), .net(N1311), .FEN(FEN[544]), .op(N1311_t2) );
fim FAN_N1315_0 ( .fault(fault), .net(N1315), .FEN(FEN[545]), .op(N1315_t0) );
fim FAN_N1315_1 ( .fault(fault), .net(N1315), .FEN(FEN[546]), .op(N1315_t1) );
fim FAN_N1315_2 ( .fault(fault), .net(N1315), .FEN(FEN[547]), .op(N1315_t2) );
fim FAN_N1319_0 ( .fault(fault), .net(N1319), .FEN(FEN[548]), .op(N1319_t0) );
fim FAN_N1319_1 ( .fault(fault), .net(N1319), .FEN(FEN[549]), .op(N1319_t1) );
fim FAN_N1319_2 ( .fault(fault), .net(N1319), .FEN(FEN[550]), .op(N1319_t2) );
fim FAN_N1323_0 ( .fault(fault), .net(N1323), .FEN(FEN[551]), .op(N1323_t0) );
fim FAN_N1323_1 ( .fault(fault), .net(N1323), .FEN(FEN[552]), .op(N1323_t1) );
fim FAN_N1323_2 ( .fault(fault), .net(N1323), .FEN(FEN[553]), .op(N1323_t2) );
fim FAN_N1327_0 ( .fault(fault), .net(N1327), .FEN(FEN[554]), .op(N1327_t0) );
fim FAN_N1327_1 ( .fault(fault), .net(N1327), .FEN(FEN[555]), .op(N1327_t1) );
fim FAN_N1327_2 ( .fault(fault), .net(N1327), .FEN(FEN[556]), .op(N1327_t2) );
fim FAN_N1331_0 ( .fault(fault), .net(N1331), .FEN(FEN[557]), .op(N1331_t0) );
fim FAN_N1331_1 ( .fault(fault), .net(N1331), .FEN(FEN[558]), .op(N1331_t1) );
fim FAN_N1331_2 ( .fault(fault), .net(N1331), .FEN(FEN[559]), .op(N1331_t2) );
fim FAN_N1335_0 ( .fault(fault), .net(N1335), .FEN(FEN[560]), .op(N1335_t0) );
fim FAN_N1335_1 ( .fault(fault), .net(N1335), .FEN(FEN[561]), .op(N1335_t1) );
fim FAN_N1335_2 ( .fault(fault), .net(N1335), .FEN(FEN[562]), .op(N1335_t2) );
fim FAN_N1339_0 ( .fault(fault), .net(N1339), .FEN(FEN[563]), .op(N1339_t0) );
fim FAN_N1339_1 ( .fault(fault), .net(N1339), .FEN(FEN[564]), .op(N1339_t1) );
fim FAN_N1339_2 ( .fault(fault), .net(N1339), .FEN(FEN[565]), .op(N1339_t2) );
fim FAN_N1343_0 ( .fault(fault), .net(N1343), .FEN(FEN[566]), .op(N1343_t0) );
fim FAN_N1343_1 ( .fault(fault), .net(N1343), .FEN(FEN[567]), .op(N1343_t1) );
fim FAN_N1343_2 ( .fault(fault), .net(N1343), .FEN(FEN[568]), .op(N1343_t2) );
fim FAN_N1347_0 ( .fault(fault), .net(N1347), .FEN(FEN[569]), .op(N1347_t0) );
fim FAN_N1347_1 ( .fault(fault), .net(N1347), .FEN(FEN[570]), .op(N1347_t1) );
fim FAN_N1347_2 ( .fault(fault), .net(N1347), .FEN(FEN[571]), .op(N1347_t2) );
fim FAN_N1351_0 ( .fault(fault), .net(N1351), .FEN(FEN[572]), .op(N1351_t0) );
fim FAN_N1351_1 ( .fault(fault), .net(N1351), .FEN(FEN[573]), .op(N1351_t1) );
fim FAN_N1351_2 ( .fault(fault), .net(N1351), .FEN(FEN[574]), .op(N1351_t2) );
fim FAN_N1355_0 ( .fault(fault), .net(N1355), .FEN(FEN[575]), .op(N1355_t0) );
fim FAN_N1355_1 ( .fault(fault), .net(N1355), .FEN(FEN[576]), .op(N1355_t1) );
fim FAN_N1355_2 ( .fault(fault), .net(N1355), .FEN(FEN[577]), .op(N1355_t2) );
fim FAN_N1359_0 ( .fault(fault), .net(N1359), .FEN(FEN[578]), .op(N1359_t0) );
fim FAN_N1359_1 ( .fault(fault), .net(N1359), .FEN(FEN[579]), .op(N1359_t1) );
fim FAN_N1359_2 ( .fault(fault), .net(N1359), .FEN(FEN[580]), .op(N1359_t2) );
fim FAN_N1363_0 ( .fault(fault), .net(N1363), .FEN(FEN[581]), .op(N1363_t0) );
fim FAN_N1363_1 ( .fault(fault), .net(N1363), .FEN(FEN[582]), .op(N1363_t1) );
fim FAN_N1363_2 ( .fault(fault), .net(N1363), .FEN(FEN[583]), .op(N1363_t2) );
fim FAN_N1367_0 ( .fault(fault), .net(N1367), .FEN(FEN[584]), .op(N1367_t0) );
fim FAN_N1367_1 ( .fault(fault), .net(N1367), .FEN(FEN[585]), .op(N1367_t1) );
fim FAN_N1367_2 ( .fault(fault), .net(N1367), .FEN(FEN[586]), .op(N1367_t2) );
fim FAN_N1401_0 ( .fault(fault), .net(N1401), .FEN(FEN[587]), .op(N1401_t0) );
fim FAN_N1401_1 ( .fault(fault), .net(N1401), .FEN(FEN[588]), .op(N1401_t1) );
fim FAN_N546_0 ( .fault(fault), .net(N546), .FEN(FEN[589]), .op(N546_t0) );
fim FAN_N546_1 ( .fault(fault), .net(N546), .FEN(FEN[590]), .op(N546_t1) );
fim FAN_N1404_0 ( .fault(fault), .net(N1404), .FEN(FEN[591]), .op(N1404_t0) );
fim FAN_N1404_1 ( .fault(fault), .net(N1404), .FEN(FEN[592]), .op(N1404_t1) );
fim FAN_N594_0 ( .fault(fault), .net(N594), .FEN(FEN[593]), .op(N594_t0) );
fim FAN_N594_1 ( .fault(fault), .net(N594), .FEN(FEN[594]), .op(N594_t1) );
fim FAN_N1407_0 ( .fault(fault), .net(N1407), .FEN(FEN[595]), .op(N1407_t0) );
fim FAN_N1407_1 ( .fault(fault), .net(N1407), .FEN(FEN[596]), .op(N1407_t1) );
fim FAN_N642_0 ( .fault(fault), .net(N642), .FEN(FEN[597]), .op(N642_t0) );
fim FAN_N642_1 ( .fault(fault), .net(N642), .FEN(FEN[598]), .op(N642_t1) );
fim FAN_N1410_0 ( .fault(fault), .net(N1410), .FEN(FEN[599]), .op(N1410_t0) );
fim FAN_N1410_1 ( .fault(fault), .net(N1410), .FEN(FEN[600]), .op(N1410_t1) );
fim FAN_N690_0 ( .fault(fault), .net(N690), .FEN(FEN[601]), .op(N690_t0) );
fim FAN_N690_1 ( .fault(fault), .net(N690), .FEN(FEN[602]), .op(N690_t1) );
fim FAN_N1413_0 ( .fault(fault), .net(N1413), .FEN(FEN[603]), .op(N1413_t0) );
fim FAN_N1413_1 ( .fault(fault), .net(N1413), .FEN(FEN[604]), .op(N1413_t1) );
fim FAN_N738_0 ( .fault(fault), .net(N738), .FEN(FEN[605]), .op(N738_t0) );
fim FAN_N738_1 ( .fault(fault), .net(N738), .FEN(FEN[606]), .op(N738_t1) );
fim FAN_N1416_0 ( .fault(fault), .net(N1416), .FEN(FEN[607]), .op(N1416_t0) );
fim FAN_N1416_1 ( .fault(fault), .net(N1416), .FEN(FEN[608]), .op(N1416_t1) );
fim FAN_N786_0 ( .fault(fault), .net(N786), .FEN(FEN[609]), .op(N786_t0) );
fim FAN_N786_1 ( .fault(fault), .net(N786), .FEN(FEN[610]), .op(N786_t1) );
fim FAN_N1419_0 ( .fault(fault), .net(N1419), .FEN(FEN[611]), .op(N1419_t0) );
fim FAN_N1419_1 ( .fault(fault), .net(N1419), .FEN(FEN[612]), .op(N1419_t1) );
fim FAN_N834_0 ( .fault(fault), .net(N834), .FEN(FEN[613]), .op(N834_t0) );
fim FAN_N834_1 ( .fault(fault), .net(N834), .FEN(FEN[614]), .op(N834_t1) );
fim FAN_N1422_0 ( .fault(fault), .net(N1422), .FEN(FEN[615]), .op(N1422_t0) );
fim FAN_N1422_1 ( .fault(fault), .net(N1422), .FEN(FEN[616]), .op(N1422_t1) );
fim FAN_N882_0 ( .fault(fault), .net(N882), .FEN(FEN[617]), .op(N882_t0) );
fim FAN_N882_1 ( .fault(fault), .net(N882), .FEN(FEN[618]), .op(N882_t1) );
fim FAN_N1425_0 ( .fault(fault), .net(N1425), .FEN(FEN[619]), .op(N1425_t0) );
fim FAN_N1425_1 ( .fault(fault), .net(N1425), .FEN(FEN[620]), .op(N1425_t1) );
fim FAN_N930_0 ( .fault(fault), .net(N930), .FEN(FEN[621]), .op(N930_t0) );
fim FAN_N930_1 ( .fault(fault), .net(N930), .FEN(FEN[622]), .op(N930_t1) );
fim FAN_N1428_0 ( .fault(fault), .net(N1428), .FEN(FEN[623]), .op(N1428_t0) );
fim FAN_N1428_1 ( .fault(fault), .net(N1428), .FEN(FEN[624]), .op(N1428_t1) );
fim FAN_N978_0 ( .fault(fault), .net(N978), .FEN(FEN[625]), .op(N978_t0) );
fim FAN_N978_1 ( .fault(fault), .net(N978), .FEN(FEN[626]), .op(N978_t1) );
fim FAN_N1431_0 ( .fault(fault), .net(N1431), .FEN(FEN[627]), .op(N1431_t0) );
fim FAN_N1431_1 ( .fault(fault), .net(N1431), .FEN(FEN[628]), .op(N1431_t1) );
fim FAN_N1026_0 ( .fault(fault), .net(N1026), .FEN(FEN[629]), .op(N1026_t0) );
fim FAN_N1026_1 ( .fault(fault), .net(N1026), .FEN(FEN[630]), .op(N1026_t1) );
fim FAN_N1434_0 ( .fault(fault), .net(N1434), .FEN(FEN[631]), .op(N1434_t0) );
fim FAN_N1434_1 ( .fault(fault), .net(N1434), .FEN(FEN[632]), .op(N1434_t1) );
fim FAN_N1074_0 ( .fault(fault), .net(N1074), .FEN(FEN[633]), .op(N1074_t0) );
fim FAN_N1074_1 ( .fault(fault), .net(N1074), .FEN(FEN[634]), .op(N1074_t1) );
fim FAN_N1437_0 ( .fault(fault), .net(N1437), .FEN(FEN[635]), .op(N1437_t0) );
fim FAN_N1437_1 ( .fault(fault), .net(N1437), .FEN(FEN[636]), .op(N1437_t1) );
fim FAN_N1122_0 ( .fault(fault), .net(N1122), .FEN(FEN[637]), .op(N1122_t0) );
fim FAN_N1122_1 ( .fault(fault), .net(N1122), .FEN(FEN[638]), .op(N1122_t1) );
fim FAN_N1440_0 ( .fault(fault), .net(N1440), .FEN(FEN[639]), .op(N1440_t0) );
fim FAN_N1440_1 ( .fault(fault), .net(N1440), .FEN(FEN[640]), .op(N1440_t1) );
fim FAN_N1170_0 ( .fault(fault), .net(N1170), .FEN(FEN[641]), .op(N1170_t0) );
fim FAN_N1170_1 ( .fault(fault), .net(N1170), .FEN(FEN[642]), .op(N1170_t1) );
fim FAN_N1443_0 ( .fault(fault), .net(N1443), .FEN(FEN[643]), .op(N1443_t0) );
fim FAN_N1443_1 ( .fault(fault), .net(N1443), .FEN(FEN[644]), .op(N1443_t1) );
fim FAN_N1218_0 ( .fault(fault), .net(N1218), .FEN(FEN[645]), .op(N1218_t0) );
fim FAN_N1218_1 ( .fault(fault), .net(N1218), .FEN(FEN[646]), .op(N1218_t1) );
fim FAN_N1446_0 ( .fault(fault), .net(N1446), .FEN(FEN[647]), .op(N1446_t0) );
fim FAN_N1446_1 ( .fault(fault), .net(N1446), .FEN(FEN[648]), .op(N1446_t1) );
fim FAN_N1446_2 ( .fault(fault), .net(N1446), .FEN(FEN[649]), .op(N1446_t2) );
fim FAN_N1450_0 ( .fault(fault), .net(N1450), .FEN(FEN[650]), .op(N1450_t0) );
fim FAN_N1450_1 ( .fault(fault), .net(N1450), .FEN(FEN[651]), .op(N1450_t1) );
fim FAN_N1450_2 ( .fault(fault), .net(N1450), .FEN(FEN[652]), .op(N1450_t2) );
fim FAN_N1454_0 ( .fault(fault), .net(N1454), .FEN(FEN[653]), .op(N1454_t0) );
fim FAN_N1454_1 ( .fault(fault), .net(N1454), .FEN(FEN[654]), .op(N1454_t1) );
fim FAN_N1454_2 ( .fault(fault), .net(N1454), .FEN(FEN[655]), .op(N1454_t2) );
fim FAN_N1458_0 ( .fault(fault), .net(N1458), .FEN(FEN[656]), .op(N1458_t0) );
fim FAN_N1458_1 ( .fault(fault), .net(N1458), .FEN(FEN[657]), .op(N1458_t1) );
fim FAN_N1458_2 ( .fault(fault), .net(N1458), .FEN(FEN[658]), .op(N1458_t2) );
fim FAN_N1462_0 ( .fault(fault), .net(N1462), .FEN(FEN[659]), .op(N1462_t0) );
fim FAN_N1462_1 ( .fault(fault), .net(N1462), .FEN(FEN[660]), .op(N1462_t1) );
fim FAN_N1462_2 ( .fault(fault), .net(N1462), .FEN(FEN[661]), .op(N1462_t2) );
fim FAN_N1466_0 ( .fault(fault), .net(N1466), .FEN(FEN[662]), .op(N1466_t0) );
fim FAN_N1466_1 ( .fault(fault), .net(N1466), .FEN(FEN[663]), .op(N1466_t1) );
fim FAN_N1466_2 ( .fault(fault), .net(N1466), .FEN(FEN[664]), .op(N1466_t2) );
fim FAN_N1470_0 ( .fault(fault), .net(N1470), .FEN(FEN[665]), .op(N1470_t0) );
fim FAN_N1470_1 ( .fault(fault), .net(N1470), .FEN(FEN[666]), .op(N1470_t1) );
fim FAN_N1470_2 ( .fault(fault), .net(N1470), .FEN(FEN[667]), .op(N1470_t2) );
fim FAN_N1474_0 ( .fault(fault), .net(N1474), .FEN(FEN[668]), .op(N1474_t0) );
fim FAN_N1474_1 ( .fault(fault), .net(N1474), .FEN(FEN[669]), .op(N1474_t1) );
fim FAN_N1474_2 ( .fault(fault), .net(N1474), .FEN(FEN[670]), .op(N1474_t2) );
fim FAN_N1478_0 ( .fault(fault), .net(N1478), .FEN(FEN[671]), .op(N1478_t0) );
fim FAN_N1478_1 ( .fault(fault), .net(N1478), .FEN(FEN[672]), .op(N1478_t1) );
fim FAN_N1478_2 ( .fault(fault), .net(N1478), .FEN(FEN[673]), .op(N1478_t2) );
fim FAN_N1482_0 ( .fault(fault), .net(N1482), .FEN(FEN[674]), .op(N1482_t0) );
fim FAN_N1482_1 ( .fault(fault), .net(N1482), .FEN(FEN[675]), .op(N1482_t1) );
fim FAN_N1482_2 ( .fault(fault), .net(N1482), .FEN(FEN[676]), .op(N1482_t2) );
fim FAN_N1486_0 ( .fault(fault), .net(N1486), .FEN(FEN[677]), .op(N1486_t0) );
fim FAN_N1486_1 ( .fault(fault), .net(N1486), .FEN(FEN[678]), .op(N1486_t1) );
fim FAN_N1486_2 ( .fault(fault), .net(N1486), .FEN(FEN[679]), .op(N1486_t2) );
fim FAN_N1490_0 ( .fault(fault), .net(N1490), .FEN(FEN[680]), .op(N1490_t0) );
fim FAN_N1490_1 ( .fault(fault), .net(N1490), .FEN(FEN[681]), .op(N1490_t1) );
fim FAN_N1490_2 ( .fault(fault), .net(N1490), .FEN(FEN[682]), .op(N1490_t2) );
fim FAN_N1494_0 ( .fault(fault), .net(N1494), .FEN(FEN[683]), .op(N1494_t0) );
fim FAN_N1494_1 ( .fault(fault), .net(N1494), .FEN(FEN[684]), .op(N1494_t1) );
fim FAN_N1494_2 ( .fault(fault), .net(N1494), .FEN(FEN[685]), .op(N1494_t2) );
fim FAN_N1498_0 ( .fault(fault), .net(N1498), .FEN(FEN[686]), .op(N1498_t0) );
fim FAN_N1498_1 ( .fault(fault), .net(N1498), .FEN(FEN[687]), .op(N1498_t1) );
fim FAN_N1498_2 ( .fault(fault), .net(N1498), .FEN(FEN[688]), .op(N1498_t2) );
fim FAN_N1502_0 ( .fault(fault), .net(N1502), .FEN(FEN[689]), .op(N1502_t0) );
fim FAN_N1502_1 ( .fault(fault), .net(N1502), .FEN(FEN[690]), .op(N1502_t1) );
fim FAN_N1502_2 ( .fault(fault), .net(N1502), .FEN(FEN[691]), .op(N1502_t2) );
fim FAN_N1266_0 ( .fault(fault), .net(N1266), .FEN(FEN[692]), .op(N1266_t0) );
fim FAN_N1266_1 ( .fault(fault), .net(N1266), .FEN(FEN[693]), .op(N1266_t1) );
fim FAN_N1578_0 ( .fault(fault), .net(N1578), .FEN(FEN[694]), .op(N1578_t0) );
fim FAN_N1578_1 ( .fault(fault), .net(N1578), .FEN(FEN[695]), .op(N1578_t1) );
fim FAN_N1582_0 ( .fault(fault), .net(N1582), .FEN(FEN[696]), .op(N1582_t0) );
fim FAN_N1582_1 ( .fault(fault), .net(N1582), .FEN(FEN[697]), .op(N1582_t1) );
fim FAN_N1508_0 ( .fault(fault), .net(N1508), .FEN(FEN[698]), .op(N1508_t0) );
fim FAN_N1508_1 ( .fault(fault), .net(N1508), .FEN(FEN[699]), .op(N1508_t1) );
fim FAN_N1585_0 ( .fault(fault), .net(N1585), .FEN(FEN[700]), .op(N1585_t0) );
fim FAN_N1585_1 ( .fault(fault), .net(N1585), .FEN(FEN[701]), .op(N1585_t1) );
fim FAN_N1513_0 ( .fault(fault), .net(N1513), .FEN(FEN[702]), .op(N1513_t0) );
fim FAN_N1513_1 ( .fault(fault), .net(N1513), .FEN(FEN[703]), .op(N1513_t1) );
fim FAN_N1588_0 ( .fault(fault), .net(N1588), .FEN(FEN[704]), .op(N1588_t0) );
fim FAN_N1588_1 ( .fault(fault), .net(N1588), .FEN(FEN[705]), .op(N1588_t1) );
fim FAN_N1518_0 ( .fault(fault), .net(N1518), .FEN(FEN[706]), .op(N1518_t0) );
fim FAN_N1518_1 ( .fault(fault), .net(N1518), .FEN(FEN[707]), .op(N1518_t1) );
fim FAN_N1591_0 ( .fault(fault), .net(N1591), .FEN(FEN[708]), .op(N1591_t0) );
fim FAN_N1591_1 ( .fault(fault), .net(N1591), .FEN(FEN[709]), .op(N1591_t1) );
fim FAN_N1523_0 ( .fault(fault), .net(N1523), .FEN(FEN[710]), .op(N1523_t0) );
fim FAN_N1523_1 ( .fault(fault), .net(N1523), .FEN(FEN[711]), .op(N1523_t1) );
fim FAN_N1594_0 ( .fault(fault), .net(N1594), .FEN(FEN[712]), .op(N1594_t0) );
fim FAN_N1594_1 ( .fault(fault), .net(N1594), .FEN(FEN[713]), .op(N1594_t1) );
fim FAN_N1528_0 ( .fault(fault), .net(N1528), .FEN(FEN[714]), .op(N1528_t0) );
fim FAN_N1528_1 ( .fault(fault), .net(N1528), .FEN(FEN[715]), .op(N1528_t1) );
fim FAN_N1597_0 ( .fault(fault), .net(N1597), .FEN(FEN[716]), .op(N1597_t0) );
fim FAN_N1597_1 ( .fault(fault), .net(N1597), .FEN(FEN[717]), .op(N1597_t1) );
fim FAN_N1533_0 ( .fault(fault), .net(N1533), .FEN(FEN[718]), .op(N1533_t0) );
fim FAN_N1533_1 ( .fault(fault), .net(N1533), .FEN(FEN[719]), .op(N1533_t1) );
fim FAN_N1600_0 ( .fault(fault), .net(N1600), .FEN(FEN[720]), .op(N1600_t0) );
fim FAN_N1600_1 ( .fault(fault), .net(N1600), .FEN(FEN[721]), .op(N1600_t1) );
fim FAN_N1538_0 ( .fault(fault), .net(N1538), .FEN(FEN[722]), .op(N1538_t0) );
fim FAN_N1538_1 ( .fault(fault), .net(N1538), .FEN(FEN[723]), .op(N1538_t1) );
fim FAN_N1603_0 ( .fault(fault), .net(N1603), .FEN(FEN[724]), .op(N1603_t0) );
fim FAN_N1603_1 ( .fault(fault), .net(N1603), .FEN(FEN[725]), .op(N1603_t1) );
fim FAN_N1543_0 ( .fault(fault), .net(N1543), .FEN(FEN[726]), .op(N1543_t0) );
fim FAN_N1543_1 ( .fault(fault), .net(N1543), .FEN(FEN[727]), .op(N1543_t1) );
fim FAN_N1606_0 ( .fault(fault), .net(N1606), .FEN(FEN[728]), .op(N1606_t0) );
fim FAN_N1606_1 ( .fault(fault), .net(N1606), .FEN(FEN[729]), .op(N1606_t1) );
fim FAN_N1548_0 ( .fault(fault), .net(N1548), .FEN(FEN[730]), .op(N1548_t0) );
fim FAN_N1548_1 ( .fault(fault), .net(N1548), .FEN(FEN[731]), .op(N1548_t1) );
fim FAN_N1609_0 ( .fault(fault), .net(N1609), .FEN(FEN[732]), .op(N1609_t0) );
fim FAN_N1609_1 ( .fault(fault), .net(N1609), .FEN(FEN[733]), .op(N1609_t1) );
fim FAN_N1553_0 ( .fault(fault), .net(N1553), .FEN(FEN[734]), .op(N1553_t0) );
fim FAN_N1553_1 ( .fault(fault), .net(N1553), .FEN(FEN[735]), .op(N1553_t1) );
fim FAN_N1612_0 ( .fault(fault), .net(N1612), .FEN(FEN[736]), .op(N1612_t0) );
fim FAN_N1612_1 ( .fault(fault), .net(N1612), .FEN(FEN[737]), .op(N1612_t1) );
fim FAN_N1558_0 ( .fault(fault), .net(N1558), .FEN(FEN[738]), .op(N1558_t0) );
fim FAN_N1558_1 ( .fault(fault), .net(N1558), .FEN(FEN[739]), .op(N1558_t1) );
fim FAN_N1615_0 ( .fault(fault), .net(N1615), .FEN(FEN[740]), .op(N1615_t0) );
fim FAN_N1615_1 ( .fault(fault), .net(N1615), .FEN(FEN[741]), .op(N1615_t1) );
fim FAN_N1563_0 ( .fault(fault), .net(N1563), .FEN(FEN[742]), .op(N1563_t0) );
fim FAN_N1563_1 ( .fault(fault), .net(N1563), .FEN(FEN[743]), .op(N1563_t1) );
fim FAN_N1618_0 ( .fault(fault), .net(N1618), .FEN(FEN[744]), .op(N1618_t0) );
fim FAN_N1618_1 ( .fault(fault), .net(N1618), .FEN(FEN[745]), .op(N1618_t1) );
fim FAN_N1568_0 ( .fault(fault), .net(N1568), .FEN(FEN[746]), .op(N1568_t0) );
fim FAN_N1568_1 ( .fault(fault), .net(N1568), .FEN(FEN[747]), .op(N1568_t1) );
fim FAN_N1621_0 ( .fault(fault), .net(N1621), .FEN(FEN[748]), .op(N1621_t0) );
fim FAN_N1621_1 ( .fault(fault), .net(N1621), .FEN(FEN[749]), .op(N1621_t1) );
fim FAN_N1573_0 ( .fault(fault), .net(N1573), .FEN(FEN[750]), .op(N1573_t0) );
fim FAN_N1573_1 ( .fault(fault), .net(N1573), .FEN(FEN[751]), .op(N1573_t1) );
fim FAN_N1624_0 ( .fault(fault), .net(N1624), .FEN(FEN[752]), .op(N1624_t0) );
fim FAN_N1624_1 ( .fault(fault), .net(N1624), .FEN(FEN[753]), .op(N1624_t1) );
fim FAN_N1624_2 ( .fault(fault), .net(N1624), .FEN(FEN[754]), .op(N1624_t2) );
fim FAN_N1628_0 ( .fault(fault), .net(N1628), .FEN(FEN[755]), .op(N1628_t0) );
fim FAN_N1628_1 ( .fault(fault), .net(N1628), .FEN(FEN[756]), .op(N1628_t1) );
fim FAN_N1628_2 ( .fault(fault), .net(N1628), .FEN(FEN[757]), .op(N1628_t2) );
fim FAN_N1632_0 ( .fault(fault), .net(N1632), .FEN(FEN[758]), .op(N1632_t0) );
fim FAN_N1632_1 ( .fault(fault), .net(N1632), .FEN(FEN[759]), .op(N1632_t1) );
fim FAN_N1632_2 ( .fault(fault), .net(N1632), .FEN(FEN[760]), .op(N1632_t2) );
fim FAN_N1636_0 ( .fault(fault), .net(N1636), .FEN(FEN[761]), .op(N1636_t0) );
fim FAN_N1636_1 ( .fault(fault), .net(N1636), .FEN(FEN[762]), .op(N1636_t1) );
fim FAN_N1636_2 ( .fault(fault), .net(N1636), .FEN(FEN[763]), .op(N1636_t2) );
fim FAN_N1640_0 ( .fault(fault), .net(N1640), .FEN(FEN[764]), .op(N1640_t0) );
fim FAN_N1640_1 ( .fault(fault), .net(N1640), .FEN(FEN[765]), .op(N1640_t1) );
fim FAN_N1640_2 ( .fault(fault), .net(N1640), .FEN(FEN[766]), .op(N1640_t2) );
fim FAN_N1644_0 ( .fault(fault), .net(N1644), .FEN(FEN[767]), .op(N1644_t0) );
fim FAN_N1644_1 ( .fault(fault), .net(N1644), .FEN(FEN[768]), .op(N1644_t1) );
fim FAN_N1644_2 ( .fault(fault), .net(N1644), .FEN(FEN[769]), .op(N1644_t2) );
fim FAN_N1648_0 ( .fault(fault), .net(N1648), .FEN(FEN[770]), .op(N1648_t0) );
fim FAN_N1648_1 ( .fault(fault), .net(N1648), .FEN(FEN[771]), .op(N1648_t1) );
fim FAN_N1648_2 ( .fault(fault), .net(N1648), .FEN(FEN[772]), .op(N1648_t2) );
fim FAN_N1652_0 ( .fault(fault), .net(N1652), .FEN(FEN[773]), .op(N1652_t0) );
fim FAN_N1652_1 ( .fault(fault), .net(N1652), .FEN(FEN[774]), .op(N1652_t1) );
fim FAN_N1652_2 ( .fault(fault), .net(N1652), .FEN(FEN[775]), .op(N1652_t2) );
fim FAN_N1656_0 ( .fault(fault), .net(N1656), .FEN(FEN[776]), .op(N1656_t0) );
fim FAN_N1656_1 ( .fault(fault), .net(N1656), .FEN(FEN[777]), .op(N1656_t1) );
fim FAN_N1656_2 ( .fault(fault), .net(N1656), .FEN(FEN[778]), .op(N1656_t2) );
fim FAN_N1660_0 ( .fault(fault), .net(N1660), .FEN(FEN[779]), .op(N1660_t0) );
fim FAN_N1660_1 ( .fault(fault), .net(N1660), .FEN(FEN[780]), .op(N1660_t1) );
fim FAN_N1660_2 ( .fault(fault), .net(N1660), .FEN(FEN[781]), .op(N1660_t2) );
fim FAN_N1664_0 ( .fault(fault), .net(N1664), .FEN(FEN[782]), .op(N1664_t0) );
fim FAN_N1664_1 ( .fault(fault), .net(N1664), .FEN(FEN[783]), .op(N1664_t1) );
fim FAN_N1664_2 ( .fault(fault), .net(N1664), .FEN(FEN[784]), .op(N1664_t2) );
fim FAN_N1668_0 ( .fault(fault), .net(N1668), .FEN(FEN[785]), .op(N1668_t0) );
fim FAN_N1668_1 ( .fault(fault), .net(N1668), .FEN(FEN[786]), .op(N1668_t1) );
fim FAN_N1668_2 ( .fault(fault), .net(N1668), .FEN(FEN[787]), .op(N1668_t2) );
fim FAN_N1672_0 ( .fault(fault), .net(N1672), .FEN(FEN[788]), .op(N1672_t0) );
fim FAN_N1672_1 ( .fault(fault), .net(N1672), .FEN(FEN[789]), .op(N1672_t1) );
fim FAN_N1672_2 ( .fault(fault), .net(N1672), .FEN(FEN[790]), .op(N1672_t2) );
fim FAN_N1676_0 ( .fault(fault), .net(N1676), .FEN(FEN[791]), .op(N1676_t0) );
fim FAN_N1676_1 ( .fault(fault), .net(N1676), .FEN(FEN[792]), .op(N1676_t1) );
fim FAN_N1676_2 ( .fault(fault), .net(N1676), .FEN(FEN[793]), .op(N1676_t2) );
fim FAN_N1680_0 ( .fault(fault), .net(N1680), .FEN(FEN[794]), .op(N1680_t0) );
fim FAN_N1680_1 ( .fault(fault), .net(N1680), .FEN(FEN[795]), .op(N1680_t1) );
fim FAN_N1680_2 ( .fault(fault), .net(N1680), .FEN(FEN[796]), .op(N1680_t2) );
fim FAN_N1714_0 ( .fault(fault), .net(N1714), .FEN(FEN[797]), .op(N1714_t0) );
fim FAN_N1714_1 ( .fault(fault), .net(N1714), .FEN(FEN[798]), .op(N1714_t1) );
fim FAN_N1221_0 ( .fault(fault), .net(N1221), .FEN(FEN[799]), .op(N1221_t0) );
fim FAN_N1221_1 ( .fault(fault), .net(N1221), .FEN(FEN[800]), .op(N1221_t1) );
fim FAN_N1717_0 ( .fault(fault), .net(N1717), .FEN(FEN[801]), .op(N1717_t0) );
fim FAN_N1717_1 ( .fault(fault), .net(N1717), .FEN(FEN[802]), .op(N1717_t1) );
fim FAN_N549_0 ( .fault(fault), .net(N549), .FEN(FEN[803]), .op(N549_t0) );
fim FAN_N549_1 ( .fault(fault), .net(N549), .FEN(FEN[804]), .op(N549_t1) );
fim FAN_N1720_0 ( .fault(fault), .net(N1720), .FEN(FEN[805]), .op(N1720_t0) );
fim FAN_N1720_1 ( .fault(fault), .net(N1720), .FEN(FEN[806]), .op(N1720_t1) );
fim FAN_N597_0 ( .fault(fault), .net(N597), .FEN(FEN[807]), .op(N597_t0) );
fim FAN_N597_1 ( .fault(fault), .net(N597), .FEN(FEN[808]), .op(N597_t1) );
fim FAN_N1723_0 ( .fault(fault), .net(N1723), .FEN(FEN[809]), .op(N1723_t0) );
fim FAN_N1723_1 ( .fault(fault), .net(N1723), .FEN(FEN[810]), .op(N1723_t1) );
fim FAN_N645_0 ( .fault(fault), .net(N645), .FEN(FEN[811]), .op(N645_t0) );
fim FAN_N645_1 ( .fault(fault), .net(N645), .FEN(FEN[812]), .op(N645_t1) );
fim FAN_N1726_0 ( .fault(fault), .net(N1726), .FEN(FEN[813]), .op(N1726_t0) );
fim FAN_N1726_1 ( .fault(fault), .net(N1726), .FEN(FEN[814]), .op(N1726_t1) );
fim FAN_N693_0 ( .fault(fault), .net(N693), .FEN(FEN[815]), .op(N693_t0) );
fim FAN_N693_1 ( .fault(fault), .net(N693), .FEN(FEN[816]), .op(N693_t1) );
fim FAN_N1729_0 ( .fault(fault), .net(N1729), .FEN(FEN[817]), .op(N1729_t0) );
fim FAN_N1729_1 ( .fault(fault), .net(N1729), .FEN(FEN[818]), .op(N1729_t1) );
fim FAN_N741_0 ( .fault(fault), .net(N741), .FEN(FEN[819]), .op(N741_t0) );
fim FAN_N741_1 ( .fault(fault), .net(N741), .FEN(FEN[820]), .op(N741_t1) );
fim FAN_N1732_0 ( .fault(fault), .net(N1732), .FEN(FEN[821]), .op(N1732_t0) );
fim FAN_N1732_1 ( .fault(fault), .net(N1732), .FEN(FEN[822]), .op(N1732_t1) );
fim FAN_N789_0 ( .fault(fault), .net(N789), .FEN(FEN[823]), .op(N789_t0) );
fim FAN_N789_1 ( .fault(fault), .net(N789), .FEN(FEN[824]), .op(N789_t1) );
fim FAN_N1735_0 ( .fault(fault), .net(N1735), .FEN(FEN[825]), .op(N1735_t0) );
fim FAN_N1735_1 ( .fault(fault), .net(N1735), .FEN(FEN[826]), .op(N1735_t1) );
fim FAN_N837_0 ( .fault(fault), .net(N837), .FEN(FEN[827]), .op(N837_t0) );
fim FAN_N837_1 ( .fault(fault), .net(N837), .FEN(FEN[828]), .op(N837_t1) );
fim FAN_N1738_0 ( .fault(fault), .net(N1738), .FEN(FEN[829]), .op(N1738_t0) );
fim FAN_N1738_1 ( .fault(fault), .net(N1738), .FEN(FEN[830]), .op(N1738_t1) );
fim FAN_N885_0 ( .fault(fault), .net(N885), .FEN(FEN[831]), .op(N885_t0) );
fim FAN_N885_1 ( .fault(fault), .net(N885), .FEN(FEN[832]), .op(N885_t1) );
fim FAN_N1741_0 ( .fault(fault), .net(N1741), .FEN(FEN[833]), .op(N1741_t0) );
fim FAN_N1741_1 ( .fault(fault), .net(N1741), .FEN(FEN[834]), .op(N1741_t1) );
fim FAN_N933_0 ( .fault(fault), .net(N933), .FEN(FEN[835]), .op(N933_t0) );
fim FAN_N933_1 ( .fault(fault), .net(N933), .FEN(FEN[836]), .op(N933_t1) );
fim FAN_N1744_0 ( .fault(fault), .net(N1744), .FEN(FEN[837]), .op(N1744_t0) );
fim FAN_N1744_1 ( .fault(fault), .net(N1744), .FEN(FEN[838]), .op(N1744_t1) );
fim FAN_N981_0 ( .fault(fault), .net(N981), .FEN(FEN[839]), .op(N981_t0) );
fim FAN_N981_1 ( .fault(fault), .net(N981), .FEN(FEN[840]), .op(N981_t1) );
fim FAN_N1747_0 ( .fault(fault), .net(N1747), .FEN(FEN[841]), .op(N1747_t0) );
fim FAN_N1747_1 ( .fault(fault), .net(N1747), .FEN(FEN[842]), .op(N1747_t1) );
fim FAN_N1029_0 ( .fault(fault), .net(N1029), .FEN(FEN[843]), .op(N1029_t0) );
fim FAN_N1029_1 ( .fault(fault), .net(N1029), .FEN(FEN[844]), .op(N1029_t1) );
fim FAN_N1750_0 ( .fault(fault), .net(N1750), .FEN(FEN[845]), .op(N1750_t0) );
fim FAN_N1750_1 ( .fault(fault), .net(N1750), .FEN(FEN[846]), .op(N1750_t1) );
fim FAN_N1077_0 ( .fault(fault), .net(N1077), .FEN(FEN[847]), .op(N1077_t0) );
fim FAN_N1077_1 ( .fault(fault), .net(N1077), .FEN(FEN[848]), .op(N1077_t1) );
fim FAN_N1753_0 ( .fault(fault), .net(N1753), .FEN(FEN[849]), .op(N1753_t0) );
fim FAN_N1753_1 ( .fault(fault), .net(N1753), .FEN(FEN[850]), .op(N1753_t1) );
fim FAN_N1125_0 ( .fault(fault), .net(N1125), .FEN(FEN[851]), .op(N1125_t0) );
fim FAN_N1125_1 ( .fault(fault), .net(N1125), .FEN(FEN[852]), .op(N1125_t1) );
fim FAN_N1756_0 ( .fault(fault), .net(N1756), .FEN(FEN[853]), .op(N1756_t0) );
fim FAN_N1756_1 ( .fault(fault), .net(N1756), .FEN(FEN[854]), .op(N1756_t1) );
fim FAN_N1173_0 ( .fault(fault), .net(N1173), .FEN(FEN[855]), .op(N1173_t0) );
fim FAN_N1173_1 ( .fault(fault), .net(N1173), .FEN(FEN[856]), .op(N1173_t1) );
fim FAN_N1759_0 ( .fault(fault), .net(N1759), .FEN(FEN[857]), .op(N1759_t0) );
fim FAN_N1759_1 ( .fault(fault), .net(N1759), .FEN(FEN[858]), .op(N1759_t1) );
fim FAN_N1759_2 ( .fault(fault), .net(N1759), .FEN(FEN[859]), .op(N1759_t2) );
fim FAN_N1763_0 ( .fault(fault), .net(N1763), .FEN(FEN[860]), .op(N1763_t0) );
fim FAN_N1763_1 ( .fault(fault), .net(N1763), .FEN(FEN[861]), .op(N1763_t1) );
fim FAN_N1763_2 ( .fault(fault), .net(N1763), .FEN(FEN[862]), .op(N1763_t2) );
fim FAN_N1767_0 ( .fault(fault), .net(N1767), .FEN(FEN[863]), .op(N1767_t0) );
fim FAN_N1767_1 ( .fault(fault), .net(N1767), .FEN(FEN[864]), .op(N1767_t1) );
fim FAN_N1767_2 ( .fault(fault), .net(N1767), .FEN(FEN[865]), .op(N1767_t2) );
fim FAN_N1771_0 ( .fault(fault), .net(N1771), .FEN(FEN[866]), .op(N1771_t0) );
fim FAN_N1771_1 ( .fault(fault), .net(N1771), .FEN(FEN[867]), .op(N1771_t1) );
fim FAN_N1771_2 ( .fault(fault), .net(N1771), .FEN(FEN[868]), .op(N1771_t2) );
fim FAN_N1775_0 ( .fault(fault), .net(N1775), .FEN(FEN[869]), .op(N1775_t0) );
fim FAN_N1775_1 ( .fault(fault), .net(N1775), .FEN(FEN[870]), .op(N1775_t1) );
fim FAN_N1775_2 ( .fault(fault), .net(N1775), .FEN(FEN[871]), .op(N1775_t2) );
fim FAN_N1779_0 ( .fault(fault), .net(N1779), .FEN(FEN[872]), .op(N1779_t0) );
fim FAN_N1779_1 ( .fault(fault), .net(N1779), .FEN(FEN[873]), .op(N1779_t1) );
fim FAN_N1779_2 ( .fault(fault), .net(N1779), .FEN(FEN[874]), .op(N1779_t2) );
fim FAN_N1783_0 ( .fault(fault), .net(N1783), .FEN(FEN[875]), .op(N1783_t0) );
fim FAN_N1783_1 ( .fault(fault), .net(N1783), .FEN(FEN[876]), .op(N1783_t1) );
fim FAN_N1783_2 ( .fault(fault), .net(N1783), .FEN(FEN[877]), .op(N1783_t2) );
fim FAN_N1787_0 ( .fault(fault), .net(N1787), .FEN(FEN[878]), .op(N1787_t0) );
fim FAN_N1787_1 ( .fault(fault), .net(N1787), .FEN(FEN[879]), .op(N1787_t1) );
fim FAN_N1787_2 ( .fault(fault), .net(N1787), .FEN(FEN[880]), .op(N1787_t2) );
fim FAN_N1791_0 ( .fault(fault), .net(N1791), .FEN(FEN[881]), .op(N1791_t0) );
fim FAN_N1791_1 ( .fault(fault), .net(N1791), .FEN(FEN[882]), .op(N1791_t1) );
fim FAN_N1791_2 ( .fault(fault), .net(N1791), .FEN(FEN[883]), .op(N1791_t2) );
fim FAN_N1795_0 ( .fault(fault), .net(N1795), .FEN(FEN[884]), .op(N1795_t0) );
fim FAN_N1795_1 ( .fault(fault), .net(N1795), .FEN(FEN[885]), .op(N1795_t1) );
fim FAN_N1795_2 ( .fault(fault), .net(N1795), .FEN(FEN[886]), .op(N1795_t2) );
fim FAN_N1799_0 ( .fault(fault), .net(N1799), .FEN(FEN[887]), .op(N1799_t0) );
fim FAN_N1799_1 ( .fault(fault), .net(N1799), .FEN(FEN[888]), .op(N1799_t1) );
fim FAN_N1799_2 ( .fault(fault), .net(N1799), .FEN(FEN[889]), .op(N1799_t2) );
fim FAN_N1803_0 ( .fault(fault), .net(N1803), .FEN(FEN[890]), .op(N1803_t0) );
fim FAN_N1803_1 ( .fault(fault), .net(N1803), .FEN(FEN[891]), .op(N1803_t1) );
fim FAN_N1803_2 ( .fault(fault), .net(N1803), .FEN(FEN[892]), .op(N1803_t2) );
fim FAN_N1807_0 ( .fault(fault), .net(N1807), .FEN(FEN[893]), .op(N1807_t0) );
fim FAN_N1807_1 ( .fault(fault), .net(N1807), .FEN(FEN[894]), .op(N1807_t1) );
fim FAN_N1807_2 ( .fault(fault), .net(N1807), .FEN(FEN[895]), .op(N1807_t2) );
fim FAN_N1811_0 ( .fault(fault), .net(N1811), .FEN(FEN[896]), .op(N1811_t0) );
fim FAN_N1811_1 ( .fault(fault), .net(N1811), .FEN(FEN[897]), .op(N1811_t1) );
fim FAN_N1811_2 ( .fault(fault), .net(N1811), .FEN(FEN[898]), .op(N1811_t2) );
fim FAN_N1815_0 ( .fault(fault), .net(N1815), .FEN(FEN[899]), .op(N1815_t0) );
fim FAN_N1815_1 ( .fault(fault), .net(N1815), .FEN(FEN[900]), .op(N1815_t1) );
fim FAN_N1815_2 ( .fault(fault), .net(N1815), .FEN(FEN[901]), .op(N1815_t2) );
fim FAN_N1269_0 ( .fault(fault), .net(N1269), .FEN(FEN[902]), .op(N1269_t0) );
fim FAN_N1269_1 ( .fault(fault), .net(N1269), .FEN(FEN[903]), .op(N1269_t1) );
fim FAN_N1821_0 ( .fault(fault), .net(N1821), .FEN(FEN[904]), .op(N1821_t0) );
fim FAN_N1821_1 ( .fault(fault), .net(N1821), .FEN(FEN[905]), .op(N1821_t1) );
fim FAN_N1894_0 ( .fault(fault), .net(N1894), .FEN(FEN[906]), .op(N1894_t0) );
fim FAN_N1894_1 ( .fault(fault), .net(N1894), .FEN(FEN[907]), .op(N1894_t1) );
fim FAN_N1891_0 ( .fault(fault), .net(N1891), .FEN(FEN[908]), .op(N1891_t0) );
fim FAN_N1891_1 ( .fault(fault), .net(N1891), .FEN(FEN[909]), .op(N1891_t1) );
fim FAN_N1897_0 ( .fault(fault), .net(N1897), .FEN(FEN[910]), .op(N1897_t0) );
fim FAN_N1897_1 ( .fault(fault), .net(N1897), .FEN(FEN[911]), .op(N1897_t1) );
fim FAN_N1897_2 ( .fault(fault), .net(N1897), .FEN(FEN[912]), .op(N1897_t2) );
fim FAN_N1902_0 ( .fault(fault), .net(N1902), .FEN(FEN[913]), .op(N1902_t0) );
fim FAN_N1902_1 ( .fault(fault), .net(N1902), .FEN(FEN[914]), .op(N1902_t1) );
fim FAN_N1826_0 ( .fault(fault), .net(N1826), .FEN(FEN[915]), .op(N1826_t0) );
fim FAN_N1826_1 ( .fault(fault), .net(N1826), .FEN(FEN[916]), .op(N1826_t1) );
fim FAN_N1905_0 ( .fault(fault), .net(N1905), .FEN(FEN[917]), .op(N1905_t0) );
fim FAN_N1905_1 ( .fault(fault), .net(N1905), .FEN(FEN[918]), .op(N1905_t1) );
fim FAN_N1831_0 ( .fault(fault), .net(N1831), .FEN(FEN[919]), .op(N1831_t0) );
fim FAN_N1831_1 ( .fault(fault), .net(N1831), .FEN(FEN[920]), .op(N1831_t1) );
fim FAN_N1908_0 ( .fault(fault), .net(N1908), .FEN(FEN[921]), .op(N1908_t0) );
fim FAN_N1908_1 ( .fault(fault), .net(N1908), .FEN(FEN[922]), .op(N1908_t1) );
fim FAN_N1836_0 ( .fault(fault), .net(N1836), .FEN(FEN[923]), .op(N1836_t0) );
fim FAN_N1836_1 ( .fault(fault), .net(N1836), .FEN(FEN[924]), .op(N1836_t1) );
fim FAN_N1911_0 ( .fault(fault), .net(N1911), .FEN(FEN[925]), .op(N1911_t0) );
fim FAN_N1911_1 ( .fault(fault), .net(N1911), .FEN(FEN[926]), .op(N1911_t1) );
fim FAN_N1841_0 ( .fault(fault), .net(N1841), .FEN(FEN[927]), .op(N1841_t0) );
fim FAN_N1841_1 ( .fault(fault), .net(N1841), .FEN(FEN[928]), .op(N1841_t1) );
fim FAN_N1914_0 ( .fault(fault), .net(N1914), .FEN(FEN[929]), .op(N1914_t0) );
fim FAN_N1914_1 ( .fault(fault), .net(N1914), .FEN(FEN[930]), .op(N1914_t1) );
fim FAN_N1846_0 ( .fault(fault), .net(N1846), .FEN(FEN[931]), .op(N1846_t0) );
fim FAN_N1846_1 ( .fault(fault), .net(N1846), .FEN(FEN[932]), .op(N1846_t1) );
fim FAN_N1917_0 ( .fault(fault), .net(N1917), .FEN(FEN[933]), .op(N1917_t0) );
fim FAN_N1917_1 ( .fault(fault), .net(N1917), .FEN(FEN[934]), .op(N1917_t1) );
fim FAN_N1851_0 ( .fault(fault), .net(N1851), .FEN(FEN[935]), .op(N1851_t0) );
fim FAN_N1851_1 ( .fault(fault), .net(N1851), .FEN(FEN[936]), .op(N1851_t1) );
fim FAN_N1920_0 ( .fault(fault), .net(N1920), .FEN(FEN[937]), .op(N1920_t0) );
fim FAN_N1920_1 ( .fault(fault), .net(N1920), .FEN(FEN[938]), .op(N1920_t1) );
fim FAN_N1856_0 ( .fault(fault), .net(N1856), .FEN(FEN[939]), .op(N1856_t0) );
fim FAN_N1856_1 ( .fault(fault), .net(N1856), .FEN(FEN[940]), .op(N1856_t1) );
fim FAN_N1923_0 ( .fault(fault), .net(N1923), .FEN(FEN[941]), .op(N1923_t0) );
fim FAN_N1923_1 ( .fault(fault), .net(N1923), .FEN(FEN[942]), .op(N1923_t1) );
fim FAN_N1861_0 ( .fault(fault), .net(N1861), .FEN(FEN[943]), .op(N1861_t0) );
fim FAN_N1861_1 ( .fault(fault), .net(N1861), .FEN(FEN[944]), .op(N1861_t1) );
fim FAN_N1926_0 ( .fault(fault), .net(N1926), .FEN(FEN[945]), .op(N1926_t0) );
fim FAN_N1926_1 ( .fault(fault), .net(N1926), .FEN(FEN[946]), .op(N1926_t1) );
fim FAN_N1866_0 ( .fault(fault), .net(N1866), .FEN(FEN[947]), .op(N1866_t0) );
fim FAN_N1866_1 ( .fault(fault), .net(N1866), .FEN(FEN[948]), .op(N1866_t1) );
fim FAN_N1929_0 ( .fault(fault), .net(N1929), .FEN(FEN[949]), .op(N1929_t0) );
fim FAN_N1929_1 ( .fault(fault), .net(N1929), .FEN(FEN[950]), .op(N1929_t1) );
fim FAN_N1871_0 ( .fault(fault), .net(N1871), .FEN(FEN[951]), .op(N1871_t0) );
fim FAN_N1871_1 ( .fault(fault), .net(N1871), .FEN(FEN[952]), .op(N1871_t1) );
fim FAN_N1932_0 ( .fault(fault), .net(N1932), .FEN(FEN[953]), .op(N1932_t0) );
fim FAN_N1932_1 ( .fault(fault), .net(N1932), .FEN(FEN[954]), .op(N1932_t1) );
fim FAN_N1876_0 ( .fault(fault), .net(N1876), .FEN(FEN[955]), .op(N1876_t0) );
fim FAN_N1876_1 ( .fault(fault), .net(N1876), .FEN(FEN[956]), .op(N1876_t1) );
fim FAN_N1935_0 ( .fault(fault), .net(N1935), .FEN(FEN[957]), .op(N1935_t0) );
fim FAN_N1935_1 ( .fault(fault), .net(N1935), .FEN(FEN[958]), .op(N1935_t1) );
fim FAN_N1881_0 ( .fault(fault), .net(N1881), .FEN(FEN[959]), .op(N1881_t0) );
fim FAN_N1881_1 ( .fault(fault), .net(N1881), .FEN(FEN[960]), .op(N1881_t1) );
fim FAN_N1938_0 ( .fault(fault), .net(N1938), .FEN(FEN[961]), .op(N1938_t0) );
fim FAN_N1938_1 ( .fault(fault), .net(N1938), .FEN(FEN[962]), .op(N1938_t1) );
fim FAN_N1886_0 ( .fault(fault), .net(N1886), .FEN(FEN[963]), .op(N1886_t0) );
fim FAN_N1886_1 ( .fault(fault), .net(N1886), .FEN(FEN[964]), .op(N1886_t1) );
fim FAN_N1941_0 ( .fault(fault), .net(N1941), .FEN(FEN[965]), .op(N1941_t0) );
fim FAN_N1941_1 ( .fault(fault), .net(N1941), .FEN(FEN[966]), .op(N1941_t1) );
fim FAN_N1941_2 ( .fault(fault), .net(N1941), .FEN(FEN[967]), .op(N1941_t2) );
fim FAN_N1947_0 ( .fault(fault), .net(N1947), .FEN(FEN[968]), .op(N1947_t0) );
fim FAN_N1947_1 ( .fault(fault), .net(N1947), .FEN(FEN[969]), .op(N1947_t1) );
fim FAN_N1947_2 ( .fault(fault), .net(N1947), .FEN(FEN[970]), .op(N1947_t2) );
fim FAN_N1951_0 ( .fault(fault), .net(N1951), .FEN(FEN[971]), .op(N1951_t0) );
fim FAN_N1951_1 ( .fault(fault), .net(N1951), .FEN(FEN[972]), .op(N1951_t1) );
fim FAN_N1951_2 ( .fault(fault), .net(N1951), .FEN(FEN[973]), .op(N1951_t2) );
fim FAN_N1955_0 ( .fault(fault), .net(N1955), .FEN(FEN[974]), .op(N1955_t0) );
fim FAN_N1955_1 ( .fault(fault), .net(N1955), .FEN(FEN[975]), .op(N1955_t1) );
fim FAN_N1955_2 ( .fault(fault), .net(N1955), .FEN(FEN[976]), .op(N1955_t2) );
fim FAN_N1959_0 ( .fault(fault), .net(N1959), .FEN(FEN[977]), .op(N1959_t0) );
fim FAN_N1959_1 ( .fault(fault), .net(N1959), .FEN(FEN[978]), .op(N1959_t1) );
fim FAN_N1959_2 ( .fault(fault), .net(N1959), .FEN(FEN[979]), .op(N1959_t2) );
fim FAN_N1963_0 ( .fault(fault), .net(N1963), .FEN(FEN[980]), .op(N1963_t0) );
fim FAN_N1963_1 ( .fault(fault), .net(N1963), .FEN(FEN[981]), .op(N1963_t1) );
fim FAN_N1963_2 ( .fault(fault), .net(N1963), .FEN(FEN[982]), .op(N1963_t2) );
fim FAN_N1967_0 ( .fault(fault), .net(N1967), .FEN(FEN[983]), .op(N1967_t0) );
fim FAN_N1967_1 ( .fault(fault), .net(N1967), .FEN(FEN[984]), .op(N1967_t1) );
fim FAN_N1967_2 ( .fault(fault), .net(N1967), .FEN(FEN[985]), .op(N1967_t2) );
fim FAN_N1971_0 ( .fault(fault), .net(N1971), .FEN(FEN[986]), .op(N1971_t0) );
fim FAN_N1971_1 ( .fault(fault), .net(N1971), .FEN(FEN[987]), .op(N1971_t1) );
fim FAN_N1971_2 ( .fault(fault), .net(N1971), .FEN(FEN[988]), .op(N1971_t2) );
fim FAN_N1975_0 ( .fault(fault), .net(N1975), .FEN(FEN[989]), .op(N1975_t0) );
fim FAN_N1975_1 ( .fault(fault), .net(N1975), .FEN(FEN[990]), .op(N1975_t1) );
fim FAN_N1975_2 ( .fault(fault), .net(N1975), .FEN(FEN[991]), .op(N1975_t2) );
fim FAN_N1979_0 ( .fault(fault), .net(N1979), .FEN(FEN[992]), .op(N1979_t0) );
fim FAN_N1979_1 ( .fault(fault), .net(N1979), .FEN(FEN[993]), .op(N1979_t1) );
fim FAN_N1979_2 ( .fault(fault), .net(N1979), .FEN(FEN[994]), .op(N1979_t2) );
fim FAN_N1983_0 ( .fault(fault), .net(N1983), .FEN(FEN[995]), .op(N1983_t0) );
fim FAN_N1983_1 ( .fault(fault), .net(N1983), .FEN(FEN[996]), .op(N1983_t1) );
fim FAN_N1983_2 ( .fault(fault), .net(N1983), .FEN(FEN[997]), .op(N1983_t2) );
fim FAN_N1987_0 ( .fault(fault), .net(N1987), .FEN(FEN[998]), .op(N1987_t0) );
fim FAN_N1987_1 ( .fault(fault), .net(N1987), .FEN(FEN[999]), .op(N1987_t1) );
fim FAN_N1987_2 ( .fault(fault), .net(N1987), .FEN(FEN[1000]), .op(N1987_t2) );
fim FAN_N1991_0 ( .fault(fault), .net(N1991), .FEN(FEN[1001]), .op(N1991_t0) );
fim FAN_N1991_1 ( .fault(fault), .net(N1991), .FEN(FEN[1002]), .op(N1991_t1) );
fim FAN_N1991_2 ( .fault(fault), .net(N1991), .FEN(FEN[1003]), .op(N1991_t2) );
fim FAN_N1995_0 ( .fault(fault), .net(N1995), .FEN(FEN[1004]), .op(N1995_t0) );
fim FAN_N1995_1 ( .fault(fault), .net(N1995), .FEN(FEN[1005]), .op(N1995_t1) );
fim FAN_N1995_2 ( .fault(fault), .net(N1995), .FEN(FEN[1006]), .op(N1995_t2) );
fim FAN_N2001_0 ( .fault(fault), .net(N2001), .FEN(FEN[1007]), .op(N2001_t0) );
fim FAN_N2001_1 ( .fault(fault), .net(N2001), .FEN(FEN[1008]), .op(N2001_t1) );
fim FAN_N1224_0 ( .fault(fault), .net(N1224), .FEN(FEN[1009]), .op(N1224_t0) );
fim FAN_N1224_1 ( .fault(fault), .net(N1224), .FEN(FEN[1010]), .op(N1224_t1) );
fim FAN_N2030_0 ( .fault(fault), .net(N2030), .FEN(FEN[1011]), .op(N2030_t0) );
fim FAN_N2030_1 ( .fault(fault), .net(N2030), .FEN(FEN[1012]), .op(N2030_t1) );
fim FAN_N1176_0 ( .fault(fault), .net(N1176), .FEN(FEN[1013]), .op(N1176_t0) );
fim FAN_N1176_1 ( .fault(fault), .net(N1176), .FEN(FEN[1014]), .op(N1176_t1) );
fim FAN_N2033_0 ( .fault(fault), .net(N2033), .FEN(FEN[1015]), .op(N2033_t0) );
fim FAN_N2033_1 ( .fault(fault), .net(N2033), .FEN(FEN[1016]), .op(N2033_t1) );
fim FAN_N2033_2 ( .fault(fault), .net(N2033), .FEN(FEN[1017]), .op(N2033_t2) );
fim FAN_N2037_0 ( .fault(fault), .net(N2037), .FEN(FEN[1018]), .op(N2037_t0) );
fim FAN_N2037_1 ( .fault(fault), .net(N2037), .FEN(FEN[1019]), .op(N2037_t1) );
fim FAN_N552_0 ( .fault(fault), .net(N552), .FEN(FEN[1020]), .op(N552_t0) );
fim FAN_N552_1 ( .fault(fault), .net(N552), .FEN(FEN[1021]), .op(N552_t1) );
fim FAN_N2040_0 ( .fault(fault), .net(N2040), .FEN(FEN[1022]), .op(N2040_t0) );
fim FAN_N2040_1 ( .fault(fault), .net(N2040), .FEN(FEN[1023]), .op(N2040_t1) );
fim FAN_N600_0 ( .fault(fault), .net(N600), .FEN(FEN[1024]), .op(N600_t0) );
fim FAN_N600_1 ( .fault(fault), .net(N600), .FEN(FEN[1025]), .op(N600_t1) );
fim FAN_N2043_0 ( .fault(fault), .net(N2043), .FEN(FEN[1026]), .op(N2043_t0) );
fim FAN_N2043_1 ( .fault(fault), .net(N2043), .FEN(FEN[1027]), .op(N2043_t1) );
fim FAN_N648_0 ( .fault(fault), .net(N648), .FEN(FEN[1028]), .op(N648_t0) );
fim FAN_N648_1 ( .fault(fault), .net(N648), .FEN(FEN[1029]), .op(N648_t1) );
fim FAN_N2046_0 ( .fault(fault), .net(N2046), .FEN(FEN[1030]), .op(N2046_t0) );
fim FAN_N2046_1 ( .fault(fault), .net(N2046), .FEN(FEN[1031]), .op(N2046_t1) );
fim FAN_N696_0 ( .fault(fault), .net(N696), .FEN(FEN[1032]), .op(N696_t0) );
fim FAN_N696_1 ( .fault(fault), .net(N696), .FEN(FEN[1033]), .op(N696_t1) );
fim FAN_N2049_0 ( .fault(fault), .net(N2049), .FEN(FEN[1034]), .op(N2049_t0) );
fim FAN_N2049_1 ( .fault(fault), .net(N2049), .FEN(FEN[1035]), .op(N2049_t1) );
fim FAN_N744_0 ( .fault(fault), .net(N744), .FEN(FEN[1036]), .op(N744_t0) );
fim FAN_N744_1 ( .fault(fault), .net(N744), .FEN(FEN[1037]), .op(N744_t1) );
fim FAN_N2052_0 ( .fault(fault), .net(N2052), .FEN(FEN[1038]), .op(N2052_t0) );
fim FAN_N2052_1 ( .fault(fault), .net(N2052), .FEN(FEN[1039]), .op(N2052_t1) );
fim FAN_N792_0 ( .fault(fault), .net(N792), .FEN(FEN[1040]), .op(N792_t0) );
fim FAN_N792_1 ( .fault(fault), .net(N792), .FEN(FEN[1041]), .op(N792_t1) );
fim FAN_N2055_0 ( .fault(fault), .net(N2055), .FEN(FEN[1042]), .op(N2055_t0) );
fim FAN_N2055_1 ( .fault(fault), .net(N2055), .FEN(FEN[1043]), .op(N2055_t1) );
fim FAN_N840_0 ( .fault(fault), .net(N840), .FEN(FEN[1044]), .op(N840_t0) );
fim FAN_N840_1 ( .fault(fault), .net(N840), .FEN(FEN[1045]), .op(N840_t1) );
fim FAN_N2058_0 ( .fault(fault), .net(N2058), .FEN(FEN[1046]), .op(N2058_t0) );
fim FAN_N2058_1 ( .fault(fault), .net(N2058), .FEN(FEN[1047]), .op(N2058_t1) );
fim FAN_N888_0 ( .fault(fault), .net(N888), .FEN(FEN[1048]), .op(N888_t0) );
fim FAN_N888_1 ( .fault(fault), .net(N888), .FEN(FEN[1049]), .op(N888_t1) );
fim FAN_N2061_0 ( .fault(fault), .net(N2061), .FEN(FEN[1050]), .op(N2061_t0) );
fim FAN_N2061_1 ( .fault(fault), .net(N2061), .FEN(FEN[1051]), .op(N2061_t1) );
fim FAN_N936_0 ( .fault(fault), .net(N936), .FEN(FEN[1052]), .op(N936_t0) );
fim FAN_N936_1 ( .fault(fault), .net(N936), .FEN(FEN[1053]), .op(N936_t1) );
fim FAN_N2064_0 ( .fault(fault), .net(N2064), .FEN(FEN[1054]), .op(N2064_t0) );
fim FAN_N2064_1 ( .fault(fault), .net(N2064), .FEN(FEN[1055]), .op(N2064_t1) );
fim FAN_N984_0 ( .fault(fault), .net(N984), .FEN(FEN[1056]), .op(N984_t0) );
fim FAN_N984_1 ( .fault(fault), .net(N984), .FEN(FEN[1057]), .op(N984_t1) );
fim FAN_N2067_0 ( .fault(fault), .net(N2067), .FEN(FEN[1058]), .op(N2067_t0) );
fim FAN_N2067_1 ( .fault(fault), .net(N2067), .FEN(FEN[1059]), .op(N2067_t1) );
fim FAN_N1032_0 ( .fault(fault), .net(N1032), .FEN(FEN[1060]), .op(N1032_t0) );
fim FAN_N1032_1 ( .fault(fault), .net(N1032), .FEN(FEN[1061]), .op(N1032_t1) );
fim FAN_N2070_0 ( .fault(fault), .net(N2070), .FEN(FEN[1062]), .op(N2070_t0) );
fim FAN_N2070_1 ( .fault(fault), .net(N2070), .FEN(FEN[1063]), .op(N2070_t1) );
fim FAN_N1080_0 ( .fault(fault), .net(N1080), .FEN(FEN[1064]), .op(N1080_t0) );
fim FAN_N1080_1 ( .fault(fault), .net(N1080), .FEN(FEN[1065]), .op(N1080_t1) );
fim FAN_N2073_0 ( .fault(fault), .net(N2073), .FEN(FEN[1066]), .op(N2073_t0) );
fim FAN_N2073_1 ( .fault(fault), .net(N2073), .FEN(FEN[1067]), .op(N2073_t1) );
fim FAN_N1128_0 ( .fault(fault), .net(N1128), .FEN(FEN[1068]), .op(N1128_t0) );
fim FAN_N1128_1 ( .fault(fault), .net(N1128), .FEN(FEN[1069]), .op(N1128_t1) );
fim FAN_N2076_0 ( .fault(fault), .net(N2076), .FEN(FEN[1070]), .op(N2076_t0) );
fim FAN_N2076_1 ( .fault(fault), .net(N2076), .FEN(FEN[1071]), .op(N2076_t1) );
fim FAN_N2076_2 ( .fault(fault), .net(N2076), .FEN(FEN[1072]), .op(N2076_t2) );
fim FAN_N1272_0 ( .fault(fault), .net(N1272), .FEN(FEN[1073]), .op(N1272_t0) );
fim FAN_N1272_1 ( .fault(fault), .net(N1272), .FEN(FEN[1074]), .op(N1272_t1) );
fim FAN_N2082_0 ( .fault(fault), .net(N2082), .FEN(FEN[1075]), .op(N2082_t0) );
fim FAN_N2082_1 ( .fault(fault), .net(N2082), .FEN(FEN[1076]), .op(N2082_t1) );
fim FAN_N2085_0 ( .fault(fault), .net(N2085), .FEN(FEN[1077]), .op(N2085_t0) );
fim FAN_N2085_1 ( .fault(fault), .net(N2085), .FEN(FEN[1078]), .op(N2085_t1) );
fim FAN_N2085_2 ( .fault(fault), .net(N2085), .FEN(FEN[1079]), .op(N2085_t2) );
fim FAN_N2089_0 ( .fault(fault), .net(N2089), .FEN(FEN[1080]), .op(N2089_t0) );
fim FAN_N2089_1 ( .fault(fault), .net(N2089), .FEN(FEN[1081]), .op(N2089_t1) );
fim FAN_N2089_2 ( .fault(fault), .net(N2089), .FEN(FEN[1082]), .op(N2089_t2) );
fim FAN_N2093_0 ( .fault(fault), .net(N2093), .FEN(FEN[1083]), .op(N2093_t0) );
fim FAN_N2093_1 ( .fault(fault), .net(N2093), .FEN(FEN[1084]), .op(N2093_t1) );
fim FAN_N2093_2 ( .fault(fault), .net(N2093), .FEN(FEN[1085]), .op(N2093_t2) );
fim FAN_N2097_0 ( .fault(fault), .net(N2097), .FEN(FEN[1086]), .op(N2097_t0) );
fim FAN_N2097_1 ( .fault(fault), .net(N2097), .FEN(FEN[1087]), .op(N2097_t1) );
fim FAN_N2097_2 ( .fault(fault), .net(N2097), .FEN(FEN[1088]), .op(N2097_t2) );
fim FAN_N2101_0 ( .fault(fault), .net(N2101), .FEN(FEN[1089]), .op(N2101_t0) );
fim FAN_N2101_1 ( .fault(fault), .net(N2101), .FEN(FEN[1090]), .op(N2101_t1) );
fim FAN_N2101_2 ( .fault(fault), .net(N2101), .FEN(FEN[1091]), .op(N2101_t2) );
fim FAN_N2105_0 ( .fault(fault), .net(N2105), .FEN(FEN[1092]), .op(N2105_t0) );
fim FAN_N2105_1 ( .fault(fault), .net(N2105), .FEN(FEN[1093]), .op(N2105_t1) );
fim FAN_N2105_2 ( .fault(fault), .net(N2105), .FEN(FEN[1094]), .op(N2105_t2) );
fim FAN_N2109_0 ( .fault(fault), .net(N2109), .FEN(FEN[1095]), .op(N2109_t0) );
fim FAN_N2109_1 ( .fault(fault), .net(N2109), .FEN(FEN[1096]), .op(N2109_t1) );
fim FAN_N2109_2 ( .fault(fault), .net(N2109), .FEN(FEN[1097]), .op(N2109_t2) );
fim FAN_N2113_0 ( .fault(fault), .net(N2113), .FEN(FEN[1098]), .op(N2113_t0) );
fim FAN_N2113_1 ( .fault(fault), .net(N2113), .FEN(FEN[1099]), .op(N2113_t1) );
fim FAN_N2113_2 ( .fault(fault), .net(N2113), .FEN(FEN[1100]), .op(N2113_t2) );
fim FAN_N2117_0 ( .fault(fault), .net(N2117), .FEN(FEN[1101]), .op(N2117_t0) );
fim FAN_N2117_1 ( .fault(fault), .net(N2117), .FEN(FEN[1102]), .op(N2117_t1) );
fim FAN_N2117_2 ( .fault(fault), .net(N2117), .FEN(FEN[1103]), .op(N2117_t2) );
fim FAN_N2121_0 ( .fault(fault), .net(N2121), .FEN(FEN[1104]), .op(N2121_t0) );
fim FAN_N2121_1 ( .fault(fault), .net(N2121), .FEN(FEN[1105]), .op(N2121_t1) );
fim FAN_N2121_2 ( .fault(fault), .net(N2121), .FEN(FEN[1106]), .op(N2121_t2) );
fim FAN_N2125_0 ( .fault(fault), .net(N2125), .FEN(FEN[1107]), .op(N2125_t0) );
fim FAN_N2125_1 ( .fault(fault), .net(N2125), .FEN(FEN[1108]), .op(N2125_t1) );
fim FAN_N2125_2 ( .fault(fault), .net(N2125), .FEN(FEN[1109]), .op(N2125_t2) );
fim FAN_N2129_0 ( .fault(fault), .net(N2129), .FEN(FEN[1110]), .op(N2129_t0) );
fim FAN_N2129_1 ( .fault(fault), .net(N2129), .FEN(FEN[1111]), .op(N2129_t1) );
fim FAN_N2129_2 ( .fault(fault), .net(N2129), .FEN(FEN[1112]), .op(N2129_t2) );
fim FAN_N2133_0 ( .fault(fault), .net(N2133), .FEN(FEN[1113]), .op(N2133_t0) );
fim FAN_N2133_1 ( .fault(fault), .net(N2133), .FEN(FEN[1114]), .op(N2133_t1) );
fim FAN_N2133_2 ( .fault(fault), .net(N2133), .FEN(FEN[1115]), .op(N2133_t2) );
fim FAN_N2142_0 ( .fault(fault), .net(N2142), .FEN(FEN[1116]), .op(N2142_t0) );
fim FAN_N2142_1 ( .fault(fault), .net(N2142), .FEN(FEN[1117]), .op(N2142_t1) );
fim FAN_N2139_0 ( .fault(fault), .net(N2139), .FEN(FEN[1118]), .op(N2139_t0) );
fim FAN_N2139_1 ( .fault(fault), .net(N2139), .FEN(FEN[1119]), .op(N2139_t1) );
fim FAN_N2145_0 ( .fault(fault), .net(N2145), .FEN(FEN[1120]), .op(N2145_t0) );
fim FAN_N2145_1 ( .fault(fault), .net(N2145), .FEN(FEN[1121]), .op(N2145_t1) );
fim FAN_N2145_2 ( .fault(fault), .net(N2145), .FEN(FEN[1122]), .op(N2145_t2) );
fim FAN_N2214_0 ( .fault(fault), .net(N2214), .FEN(FEN[1123]), .op(N2214_t0) );
fim FAN_N2214_1 ( .fault(fault), .net(N2214), .FEN(FEN[1124]), .op(N2214_t1) );
fim FAN_N2211_0 ( .fault(fault), .net(N2211), .FEN(FEN[1125]), .op(N2211_t0) );
fim FAN_N2211_1 ( .fault(fault), .net(N2211), .FEN(FEN[1126]), .op(N2211_t1) );
fim FAN_N2217_0 ( .fault(fault), .net(N2217), .FEN(FEN[1127]), .op(N2217_t0) );
fim FAN_N2217_1 ( .fault(fault), .net(N2217), .FEN(FEN[1128]), .op(N2217_t1) );
fim FAN_N2217_2 ( .fault(fault), .net(N2217), .FEN(FEN[1129]), .op(N2217_t2) );
fim FAN_N2224_0 ( .fault(fault), .net(N2224), .FEN(FEN[1130]), .op(N2224_t0) );
fim FAN_N2224_1 ( .fault(fault), .net(N2224), .FEN(FEN[1131]), .op(N2224_t1) );
fim FAN_N2151_0 ( .fault(fault), .net(N2151), .FEN(FEN[1132]), .op(N2151_t0) );
fim FAN_N2151_1 ( .fault(fault), .net(N2151), .FEN(FEN[1133]), .op(N2151_t1) );
fim FAN_N2227_0 ( .fault(fault), .net(N2227), .FEN(FEN[1134]), .op(N2227_t0) );
fim FAN_N2227_1 ( .fault(fault), .net(N2227), .FEN(FEN[1135]), .op(N2227_t1) );
fim FAN_N2156_0 ( .fault(fault), .net(N2156), .FEN(FEN[1136]), .op(N2156_t0) );
fim FAN_N2156_1 ( .fault(fault), .net(N2156), .FEN(FEN[1137]), .op(N2156_t1) );
fim FAN_N2230_0 ( .fault(fault), .net(N2230), .FEN(FEN[1138]), .op(N2230_t0) );
fim FAN_N2230_1 ( .fault(fault), .net(N2230), .FEN(FEN[1139]), .op(N2230_t1) );
fim FAN_N2161_0 ( .fault(fault), .net(N2161), .FEN(FEN[1140]), .op(N2161_t0) );
fim FAN_N2161_1 ( .fault(fault), .net(N2161), .FEN(FEN[1141]), .op(N2161_t1) );
fim FAN_N2233_0 ( .fault(fault), .net(N2233), .FEN(FEN[1142]), .op(N2233_t0) );
fim FAN_N2233_1 ( .fault(fault), .net(N2233), .FEN(FEN[1143]), .op(N2233_t1) );
fim FAN_N2166_0 ( .fault(fault), .net(N2166), .FEN(FEN[1144]), .op(N2166_t0) );
fim FAN_N2166_1 ( .fault(fault), .net(N2166), .FEN(FEN[1145]), .op(N2166_t1) );
fim FAN_N2236_0 ( .fault(fault), .net(N2236), .FEN(FEN[1146]), .op(N2236_t0) );
fim FAN_N2236_1 ( .fault(fault), .net(N2236), .FEN(FEN[1147]), .op(N2236_t1) );
fim FAN_N2171_0 ( .fault(fault), .net(N2171), .FEN(FEN[1148]), .op(N2171_t0) );
fim FAN_N2171_1 ( .fault(fault), .net(N2171), .FEN(FEN[1149]), .op(N2171_t1) );
fim FAN_N2239_0 ( .fault(fault), .net(N2239), .FEN(FEN[1150]), .op(N2239_t0) );
fim FAN_N2239_1 ( .fault(fault), .net(N2239), .FEN(FEN[1151]), .op(N2239_t1) );
fim FAN_N2176_0 ( .fault(fault), .net(N2176), .FEN(FEN[1152]), .op(N2176_t0) );
fim FAN_N2176_1 ( .fault(fault), .net(N2176), .FEN(FEN[1153]), .op(N2176_t1) );
fim FAN_N2242_0 ( .fault(fault), .net(N2242), .FEN(FEN[1154]), .op(N2242_t0) );
fim FAN_N2242_1 ( .fault(fault), .net(N2242), .FEN(FEN[1155]), .op(N2242_t1) );
fim FAN_N2181_0 ( .fault(fault), .net(N2181), .FEN(FEN[1156]), .op(N2181_t0) );
fim FAN_N2181_1 ( .fault(fault), .net(N2181), .FEN(FEN[1157]), .op(N2181_t1) );
fim FAN_N2245_0 ( .fault(fault), .net(N2245), .FEN(FEN[1158]), .op(N2245_t0) );
fim FAN_N2245_1 ( .fault(fault), .net(N2245), .FEN(FEN[1159]), .op(N2245_t1) );
fim FAN_N2186_0 ( .fault(fault), .net(N2186), .FEN(FEN[1160]), .op(N2186_t0) );
fim FAN_N2186_1 ( .fault(fault), .net(N2186), .FEN(FEN[1161]), .op(N2186_t1) );
fim FAN_N2248_0 ( .fault(fault), .net(N2248), .FEN(FEN[1162]), .op(N2248_t0) );
fim FAN_N2248_1 ( .fault(fault), .net(N2248), .FEN(FEN[1163]), .op(N2248_t1) );
fim FAN_N2191_0 ( .fault(fault), .net(N2191), .FEN(FEN[1164]), .op(N2191_t0) );
fim FAN_N2191_1 ( .fault(fault), .net(N2191), .FEN(FEN[1165]), .op(N2191_t1) );
fim FAN_N2251_0 ( .fault(fault), .net(N2251), .FEN(FEN[1166]), .op(N2251_t0) );
fim FAN_N2251_1 ( .fault(fault), .net(N2251), .FEN(FEN[1167]), .op(N2251_t1) );
fim FAN_N2196_0 ( .fault(fault), .net(N2196), .FEN(FEN[1168]), .op(N2196_t0) );
fim FAN_N2196_1 ( .fault(fault), .net(N2196), .FEN(FEN[1169]), .op(N2196_t1) );
fim FAN_N2254_0 ( .fault(fault), .net(N2254), .FEN(FEN[1170]), .op(N2254_t0) );
fim FAN_N2254_1 ( .fault(fault), .net(N2254), .FEN(FEN[1171]), .op(N2254_t1) );
fim FAN_N2201_0 ( .fault(fault), .net(N2201), .FEN(FEN[1172]), .op(N2201_t0) );
fim FAN_N2201_1 ( .fault(fault), .net(N2201), .FEN(FEN[1173]), .op(N2201_t1) );
fim FAN_N2257_0 ( .fault(fault), .net(N2257), .FEN(FEN[1174]), .op(N2257_t0) );
fim FAN_N2257_1 ( .fault(fault), .net(N2257), .FEN(FEN[1175]), .op(N2257_t1) );
fim FAN_N2206_0 ( .fault(fault), .net(N2206), .FEN(FEN[1176]), .op(N2206_t0) );
fim FAN_N2206_1 ( .fault(fault), .net(N2206), .FEN(FEN[1177]), .op(N2206_t1) );
fim FAN_N2260_0 ( .fault(fault), .net(N2260), .FEN(FEN[1178]), .op(N2260_t0) );
fim FAN_N2260_1 ( .fault(fault), .net(N2260), .FEN(FEN[1179]), .op(N2260_t1) );
fim FAN_N2260_2 ( .fault(fault), .net(N2260), .FEN(FEN[1180]), .op(N2260_t2) );
fim FAN_N2266_0 ( .fault(fault), .net(N2266), .FEN(FEN[1181]), .op(N2266_t0) );
fim FAN_N2266_1 ( .fault(fault), .net(N2266), .FEN(FEN[1182]), .op(N2266_t1) );
fim FAN_N1227_0 ( .fault(fault), .net(N1227), .FEN(FEN[1183]), .op(N1227_t0) );
fim FAN_N1227_1 ( .fault(fault), .net(N1227), .FEN(FEN[1184]), .op(N1227_t1) );
fim FAN_N2269_0 ( .fault(fault), .net(N2269), .FEN(FEN[1185]), .op(N2269_t0) );
fim FAN_N2269_1 ( .fault(fault), .net(N2269), .FEN(FEN[1186]), .op(N2269_t1) );
fim FAN_N2269_2 ( .fault(fault), .net(N2269), .FEN(FEN[1187]), .op(N2269_t2) );
fim FAN_N2273_0 ( .fault(fault), .net(N2273), .FEN(FEN[1188]), .op(N2273_t0) );
fim FAN_N2273_1 ( .fault(fault), .net(N2273), .FEN(FEN[1189]), .op(N2273_t1) );
fim FAN_N2273_2 ( .fault(fault), .net(N2273), .FEN(FEN[1190]), .op(N2273_t2) );
fim FAN_N2277_0 ( .fault(fault), .net(N2277), .FEN(FEN[1191]), .op(N2277_t0) );
fim FAN_N2277_1 ( .fault(fault), .net(N2277), .FEN(FEN[1192]), .op(N2277_t1) );
fim FAN_N2277_2 ( .fault(fault), .net(N2277), .FEN(FEN[1193]), .op(N2277_t2) );
fim FAN_N2281_0 ( .fault(fault), .net(N2281), .FEN(FEN[1194]), .op(N2281_t0) );
fim FAN_N2281_1 ( .fault(fault), .net(N2281), .FEN(FEN[1195]), .op(N2281_t1) );
fim FAN_N2281_2 ( .fault(fault), .net(N2281), .FEN(FEN[1196]), .op(N2281_t2) );
fim FAN_N2285_0 ( .fault(fault), .net(N2285), .FEN(FEN[1197]), .op(N2285_t0) );
fim FAN_N2285_1 ( .fault(fault), .net(N2285), .FEN(FEN[1198]), .op(N2285_t1) );
fim FAN_N2285_2 ( .fault(fault), .net(N2285), .FEN(FEN[1199]), .op(N2285_t2) );
fim FAN_N2289_0 ( .fault(fault), .net(N2289), .FEN(FEN[1200]), .op(N2289_t0) );
fim FAN_N2289_1 ( .fault(fault), .net(N2289), .FEN(FEN[1201]), .op(N2289_t1) );
fim FAN_N2289_2 ( .fault(fault), .net(N2289), .FEN(FEN[1202]), .op(N2289_t2) );
fim FAN_N2293_0 ( .fault(fault), .net(N2293), .FEN(FEN[1203]), .op(N2293_t0) );
fim FAN_N2293_1 ( .fault(fault), .net(N2293), .FEN(FEN[1204]), .op(N2293_t1) );
fim FAN_N2293_2 ( .fault(fault), .net(N2293), .FEN(FEN[1205]), .op(N2293_t2) );
fim FAN_N2297_0 ( .fault(fault), .net(N2297), .FEN(FEN[1206]), .op(N2297_t0) );
fim FAN_N2297_1 ( .fault(fault), .net(N2297), .FEN(FEN[1207]), .op(N2297_t1) );
fim FAN_N2297_2 ( .fault(fault), .net(N2297), .FEN(FEN[1208]), .op(N2297_t2) );
fim FAN_N2301_0 ( .fault(fault), .net(N2301), .FEN(FEN[1209]), .op(N2301_t0) );
fim FAN_N2301_1 ( .fault(fault), .net(N2301), .FEN(FEN[1210]), .op(N2301_t1) );
fim FAN_N2301_2 ( .fault(fault), .net(N2301), .FEN(FEN[1211]), .op(N2301_t2) );
fim FAN_N2305_0 ( .fault(fault), .net(N2305), .FEN(FEN[1212]), .op(N2305_t0) );
fim FAN_N2305_1 ( .fault(fault), .net(N2305), .FEN(FEN[1213]), .op(N2305_t1) );
fim FAN_N2305_2 ( .fault(fault), .net(N2305), .FEN(FEN[1214]), .op(N2305_t2) );
fim FAN_N2309_0 ( .fault(fault), .net(N2309), .FEN(FEN[1215]), .op(N2309_t0) );
fim FAN_N2309_1 ( .fault(fault), .net(N2309), .FEN(FEN[1216]), .op(N2309_t1) );
fim FAN_N2309_2 ( .fault(fault), .net(N2309), .FEN(FEN[1217]), .op(N2309_t2) );
fim FAN_N2313_0 ( .fault(fault), .net(N2313), .FEN(FEN[1218]), .op(N2313_t0) );
fim FAN_N2313_1 ( .fault(fault), .net(N2313), .FEN(FEN[1219]), .op(N2313_t1) );
fim FAN_N2313_2 ( .fault(fault), .net(N2313), .FEN(FEN[1220]), .op(N2313_t2) );
fim FAN_N2319_0 ( .fault(fault), .net(N2319), .FEN(FEN[1221]), .op(N2319_t0) );
fim FAN_N2319_1 ( .fault(fault), .net(N2319), .FEN(FEN[1222]), .op(N2319_t1) );
fim FAN_N1179_0 ( .fault(fault), .net(N1179), .FEN(FEN[1223]), .op(N1179_t0) );
fim FAN_N1179_1 ( .fault(fault), .net(N1179), .FEN(FEN[1224]), .op(N1179_t1) );
fim FAN_N2322_0 ( .fault(fault), .net(N2322), .FEN(FEN[1225]), .op(N2322_t0) );
fim FAN_N2322_1 ( .fault(fault), .net(N2322), .FEN(FEN[1226]), .op(N2322_t1) );
fim FAN_N2322_2 ( .fault(fault), .net(N2322), .FEN(FEN[1227]), .op(N2322_t2) );
fim FAN_N2350_0 ( .fault(fault), .net(N2350), .FEN(FEN[1228]), .op(N2350_t0) );
fim FAN_N2350_1 ( .fault(fault), .net(N2350), .FEN(FEN[1229]), .op(N2350_t1) );
fim FAN_N1131_0 ( .fault(fault), .net(N1131), .FEN(FEN[1230]), .op(N1131_t0) );
fim FAN_N1131_1 ( .fault(fault), .net(N1131), .FEN(FEN[1231]), .op(N1131_t1) );
fim FAN_N2353_0 ( .fault(fault), .net(N2353), .FEN(FEN[1232]), .op(N2353_t0) );
fim FAN_N2353_1 ( .fault(fault), .net(N2353), .FEN(FEN[1233]), .op(N2353_t1) );
fim FAN_N2353_2 ( .fault(fault), .net(N2353), .FEN(FEN[1234]), .op(N2353_t2) );
fim FAN_N1275_0 ( .fault(fault), .net(N1275), .FEN(FEN[1235]), .op(N1275_t0) );
fim FAN_N1275_1 ( .fault(fault), .net(N1275), .FEN(FEN[1236]), .op(N1275_t1) );
fim FAN_N2359_0 ( .fault(fault), .net(N2359), .FEN(FEN[1237]), .op(N2359_t0) );
fim FAN_N2359_1 ( .fault(fault), .net(N2359), .FEN(FEN[1238]), .op(N2359_t1) );
fim FAN_N2362_0 ( .fault(fault), .net(N2362), .FEN(FEN[1239]), .op(N2362_t0) );
fim FAN_N2362_1 ( .fault(fault), .net(N2362), .FEN(FEN[1240]), .op(N2362_t1) );
fim FAN_N555_0 ( .fault(fault), .net(N555), .FEN(FEN[1241]), .op(N555_t0) );
fim FAN_N555_1 ( .fault(fault), .net(N555), .FEN(FEN[1242]), .op(N555_t1) );
fim FAN_N2365_0 ( .fault(fault), .net(N2365), .FEN(FEN[1243]), .op(N2365_t0) );
fim FAN_N2365_1 ( .fault(fault), .net(N2365), .FEN(FEN[1244]), .op(N2365_t1) );
fim FAN_N603_0 ( .fault(fault), .net(N603), .FEN(FEN[1245]), .op(N603_t0) );
fim FAN_N603_1 ( .fault(fault), .net(N603), .FEN(FEN[1246]), .op(N603_t1) );
fim FAN_N2368_0 ( .fault(fault), .net(N2368), .FEN(FEN[1247]), .op(N2368_t0) );
fim FAN_N2368_1 ( .fault(fault), .net(N2368), .FEN(FEN[1248]), .op(N2368_t1) );
fim FAN_N651_0 ( .fault(fault), .net(N651), .FEN(FEN[1249]), .op(N651_t0) );
fim FAN_N651_1 ( .fault(fault), .net(N651), .FEN(FEN[1250]), .op(N651_t1) );
fim FAN_N2371_0 ( .fault(fault), .net(N2371), .FEN(FEN[1251]), .op(N2371_t0) );
fim FAN_N2371_1 ( .fault(fault), .net(N2371), .FEN(FEN[1252]), .op(N2371_t1) );
fim FAN_N699_0 ( .fault(fault), .net(N699), .FEN(FEN[1253]), .op(N699_t0) );
fim FAN_N699_1 ( .fault(fault), .net(N699), .FEN(FEN[1254]), .op(N699_t1) );
fim FAN_N2374_0 ( .fault(fault), .net(N2374), .FEN(FEN[1255]), .op(N2374_t0) );
fim FAN_N2374_1 ( .fault(fault), .net(N2374), .FEN(FEN[1256]), .op(N2374_t1) );
fim FAN_N747_0 ( .fault(fault), .net(N747), .FEN(FEN[1257]), .op(N747_t0) );
fim FAN_N747_1 ( .fault(fault), .net(N747), .FEN(FEN[1258]), .op(N747_t1) );
fim FAN_N2377_0 ( .fault(fault), .net(N2377), .FEN(FEN[1259]), .op(N2377_t0) );
fim FAN_N2377_1 ( .fault(fault), .net(N2377), .FEN(FEN[1260]), .op(N2377_t1) );
fim FAN_N795_0 ( .fault(fault), .net(N795), .FEN(FEN[1261]), .op(N795_t0) );
fim FAN_N795_1 ( .fault(fault), .net(N795), .FEN(FEN[1262]), .op(N795_t1) );
fim FAN_N2380_0 ( .fault(fault), .net(N2380), .FEN(FEN[1263]), .op(N2380_t0) );
fim FAN_N2380_1 ( .fault(fault), .net(N2380), .FEN(FEN[1264]), .op(N2380_t1) );
fim FAN_N843_0 ( .fault(fault), .net(N843), .FEN(FEN[1265]), .op(N843_t0) );
fim FAN_N843_1 ( .fault(fault), .net(N843), .FEN(FEN[1266]), .op(N843_t1) );
fim FAN_N2383_0 ( .fault(fault), .net(N2383), .FEN(FEN[1267]), .op(N2383_t0) );
fim FAN_N2383_1 ( .fault(fault), .net(N2383), .FEN(FEN[1268]), .op(N2383_t1) );
fim FAN_N891_0 ( .fault(fault), .net(N891), .FEN(FEN[1269]), .op(N891_t0) );
fim FAN_N891_1 ( .fault(fault), .net(N891), .FEN(FEN[1270]), .op(N891_t1) );
fim FAN_N2386_0 ( .fault(fault), .net(N2386), .FEN(FEN[1271]), .op(N2386_t0) );
fim FAN_N2386_1 ( .fault(fault), .net(N2386), .FEN(FEN[1272]), .op(N2386_t1) );
fim FAN_N939_0 ( .fault(fault), .net(N939), .FEN(FEN[1273]), .op(N939_t0) );
fim FAN_N939_1 ( .fault(fault), .net(N939), .FEN(FEN[1274]), .op(N939_t1) );
fim FAN_N2389_0 ( .fault(fault), .net(N2389), .FEN(FEN[1275]), .op(N2389_t0) );
fim FAN_N2389_1 ( .fault(fault), .net(N2389), .FEN(FEN[1276]), .op(N2389_t1) );
fim FAN_N987_0 ( .fault(fault), .net(N987), .FEN(FEN[1277]), .op(N987_t0) );
fim FAN_N987_1 ( .fault(fault), .net(N987), .FEN(FEN[1278]), .op(N987_t1) );
fim FAN_N2392_0 ( .fault(fault), .net(N2392), .FEN(FEN[1279]), .op(N2392_t0) );
fim FAN_N2392_1 ( .fault(fault), .net(N2392), .FEN(FEN[1280]), .op(N2392_t1) );
fim FAN_N1035_0 ( .fault(fault), .net(N1035), .FEN(FEN[1281]), .op(N1035_t0) );
fim FAN_N1035_1 ( .fault(fault), .net(N1035), .FEN(FEN[1282]), .op(N1035_t1) );
fim FAN_N2395_0 ( .fault(fault), .net(N2395), .FEN(FEN[1283]), .op(N2395_t0) );
fim FAN_N2395_1 ( .fault(fault), .net(N2395), .FEN(FEN[1284]), .op(N2395_t1) );
fim FAN_N1083_0 ( .fault(fault), .net(N1083), .FEN(FEN[1285]), .op(N1083_t0) );
fim FAN_N1083_1 ( .fault(fault), .net(N1083), .FEN(FEN[1286]), .op(N1083_t1) );
fim FAN_N2398_0 ( .fault(fault), .net(N2398), .FEN(FEN[1287]), .op(N2398_t0) );
fim FAN_N2398_1 ( .fault(fault), .net(N2398), .FEN(FEN[1288]), .op(N2398_t1) );
fim FAN_N2398_2 ( .fault(fault), .net(N2398), .FEN(FEN[1289]), .op(N2398_t2) );
fim FAN_N2407_0 ( .fault(fault), .net(N2407), .FEN(FEN[1290]), .op(N2407_t0) );
fim FAN_N2407_1 ( .fault(fault), .net(N2407), .FEN(FEN[1291]), .op(N2407_t1) );
fim FAN_N2404_0 ( .fault(fault), .net(N2404), .FEN(FEN[1292]), .op(N2404_t0) );
fim FAN_N2404_1 ( .fault(fault), .net(N2404), .FEN(FEN[1293]), .op(N2404_t1) );
fim FAN_N2410_0 ( .fault(fault), .net(N2410), .FEN(FEN[1294]), .op(N2410_t0) );
fim FAN_N2410_1 ( .fault(fault), .net(N2410), .FEN(FEN[1295]), .op(N2410_t1) );
fim FAN_N2410_2 ( .fault(fault), .net(N2410), .FEN(FEN[1296]), .op(N2410_t2) );
fim FAN_N2414_0 ( .fault(fault), .net(N2414), .FEN(FEN[1297]), .op(N2414_t0) );
fim FAN_N2414_1 ( .fault(fault), .net(N2414), .FEN(FEN[1298]), .op(N2414_t1) );
fim FAN_N2414_2 ( .fault(fault), .net(N2414), .FEN(FEN[1299]), .op(N2414_t2) );
fim FAN_N2418_0 ( .fault(fault), .net(N2418), .FEN(FEN[1300]), .op(N2418_t0) );
fim FAN_N2418_1 ( .fault(fault), .net(N2418), .FEN(FEN[1301]), .op(N2418_t1) );
fim FAN_N2418_2 ( .fault(fault), .net(N2418), .FEN(FEN[1302]), .op(N2418_t2) );
fim FAN_N2422_0 ( .fault(fault), .net(N2422), .FEN(FEN[1303]), .op(N2422_t0) );
fim FAN_N2422_1 ( .fault(fault), .net(N2422), .FEN(FEN[1304]), .op(N2422_t1) );
fim FAN_N2422_2 ( .fault(fault), .net(N2422), .FEN(FEN[1305]), .op(N2422_t2) );
fim FAN_N2426_0 ( .fault(fault), .net(N2426), .FEN(FEN[1306]), .op(N2426_t0) );
fim FAN_N2426_1 ( .fault(fault), .net(N2426), .FEN(FEN[1307]), .op(N2426_t1) );
fim FAN_N2426_2 ( .fault(fault), .net(N2426), .FEN(FEN[1308]), .op(N2426_t2) );
fim FAN_N2430_0 ( .fault(fault), .net(N2430), .FEN(FEN[1309]), .op(N2430_t0) );
fim FAN_N2430_1 ( .fault(fault), .net(N2430), .FEN(FEN[1310]), .op(N2430_t1) );
fim FAN_N2430_2 ( .fault(fault), .net(N2430), .FEN(FEN[1311]), .op(N2430_t2) );
fim FAN_N2434_0 ( .fault(fault), .net(N2434), .FEN(FEN[1312]), .op(N2434_t0) );
fim FAN_N2434_1 ( .fault(fault), .net(N2434), .FEN(FEN[1313]), .op(N2434_t1) );
fim FAN_N2434_2 ( .fault(fault), .net(N2434), .FEN(FEN[1314]), .op(N2434_t2) );
fim FAN_N2438_0 ( .fault(fault), .net(N2438), .FEN(FEN[1315]), .op(N2438_t0) );
fim FAN_N2438_1 ( .fault(fault), .net(N2438), .FEN(FEN[1316]), .op(N2438_t1) );
fim FAN_N2438_2 ( .fault(fault), .net(N2438), .FEN(FEN[1317]), .op(N2438_t2) );
fim FAN_N2442_0 ( .fault(fault), .net(N2442), .FEN(FEN[1318]), .op(N2442_t0) );
fim FAN_N2442_1 ( .fault(fault), .net(N2442), .FEN(FEN[1319]), .op(N2442_t1) );
fim FAN_N2442_2 ( .fault(fault), .net(N2442), .FEN(FEN[1320]), .op(N2442_t2) );
fim FAN_N2446_0 ( .fault(fault), .net(N2446), .FEN(FEN[1321]), .op(N2446_t0) );
fim FAN_N2446_1 ( .fault(fault), .net(N2446), .FEN(FEN[1322]), .op(N2446_t1) );
fim FAN_N2446_2 ( .fault(fault), .net(N2446), .FEN(FEN[1323]), .op(N2446_t2) );
fim FAN_N2450_0 ( .fault(fault), .net(N2450), .FEN(FEN[1324]), .op(N2450_t0) );
fim FAN_N2450_1 ( .fault(fault), .net(N2450), .FEN(FEN[1325]), .op(N2450_t1) );
fim FAN_N2450_2 ( .fault(fault), .net(N2450), .FEN(FEN[1326]), .op(N2450_t2) );
fim FAN_N2454_0 ( .fault(fault), .net(N2454), .FEN(FEN[1327]), .op(N2454_t0) );
fim FAN_N2454_1 ( .fault(fault), .net(N2454), .FEN(FEN[1328]), .op(N2454_t1) );
fim FAN_N2454_2 ( .fault(fault), .net(N2454), .FEN(FEN[1329]), .op(N2454_t2) );
fim FAN_N2458_0 ( .fault(fault), .net(N2458), .FEN(FEN[1330]), .op(N2458_t0) );
fim FAN_N2458_1 ( .fault(fault), .net(N2458), .FEN(FEN[1331]), .op(N2458_t1) );
fim FAN_N2458_2 ( .fault(fault), .net(N2458), .FEN(FEN[1332]), .op(N2458_t2) );
fim FAN_N2467_0 ( .fault(fault), .net(N2467), .FEN(FEN[1333]), .op(N2467_t0) );
fim FAN_N2467_1 ( .fault(fault), .net(N2467), .FEN(FEN[1334]), .op(N2467_t1) );
fim FAN_N2464_0 ( .fault(fault), .net(N2464), .FEN(FEN[1335]), .op(N2464_t0) );
fim FAN_N2464_1 ( .fault(fault), .net(N2464), .FEN(FEN[1336]), .op(N2464_t1) );
fim FAN_N2470_0 ( .fault(fault), .net(N2470), .FEN(FEN[1337]), .op(N2470_t0) );
fim FAN_N2470_1 ( .fault(fault), .net(N2470), .FEN(FEN[1338]), .op(N2470_t1) );
fim FAN_N2470_2 ( .fault(fault), .net(N2470), .FEN(FEN[1339]), .op(N2470_t2) );
fim FAN_N2536_0 ( .fault(fault), .net(N2536), .FEN(FEN[1340]), .op(N2536_t0) );
fim FAN_N2536_1 ( .fault(fault), .net(N2536), .FEN(FEN[1341]), .op(N2536_t1) );
fim FAN_N2533_0 ( .fault(fault), .net(N2533), .FEN(FEN[1342]), .op(N2533_t0) );
fim FAN_N2533_1 ( .fault(fault), .net(N2533), .FEN(FEN[1343]), .op(N2533_t1) );
fim FAN_N2539_0 ( .fault(fault), .net(N2539), .FEN(FEN[1344]), .op(N2539_t0) );
fim FAN_N2539_1 ( .fault(fault), .net(N2539), .FEN(FEN[1345]), .op(N2539_t1) );
fim FAN_N2539_2 ( .fault(fault), .net(N2539), .FEN(FEN[1346]), .op(N2539_t2) );
fim FAN_N2545_0 ( .fault(fault), .net(N2545), .FEN(FEN[1347]), .op(N2545_t0) );
fim FAN_N2545_1 ( .fault(fault), .net(N2545), .FEN(FEN[1348]), .op(N2545_t1) );
fim FAN_N1230_0 ( .fault(fault), .net(N1230), .FEN(FEN[1349]), .op(N1230_t0) );
fim FAN_N1230_1 ( .fault(fault), .net(N1230), .FEN(FEN[1350]), .op(N1230_t1) );
fim FAN_N2549_0 ( .fault(fault), .net(N2549), .FEN(FEN[1351]), .op(N2549_t0) );
fim FAN_N2549_1 ( .fault(fault), .net(N2549), .FEN(FEN[1352]), .op(N2549_t1) );
fim FAN_N2478_0 ( .fault(fault), .net(N2478), .FEN(FEN[1353]), .op(N2478_t0) );
fim FAN_N2478_1 ( .fault(fault), .net(N2478), .FEN(FEN[1354]), .op(N2478_t1) );
fim FAN_N2552_0 ( .fault(fault), .net(N2552), .FEN(FEN[1355]), .op(N2552_t0) );
fim FAN_N2552_1 ( .fault(fault), .net(N2552), .FEN(FEN[1356]), .op(N2552_t1) );
fim FAN_N2483_0 ( .fault(fault), .net(N2483), .FEN(FEN[1357]), .op(N2483_t0) );
fim FAN_N2483_1 ( .fault(fault), .net(N2483), .FEN(FEN[1358]), .op(N2483_t1) );
fim FAN_N2555_0 ( .fault(fault), .net(N2555), .FEN(FEN[1359]), .op(N2555_t0) );
fim FAN_N2555_1 ( .fault(fault), .net(N2555), .FEN(FEN[1360]), .op(N2555_t1) );
fim FAN_N2488_0 ( .fault(fault), .net(N2488), .FEN(FEN[1361]), .op(N2488_t0) );
fim FAN_N2488_1 ( .fault(fault), .net(N2488), .FEN(FEN[1362]), .op(N2488_t1) );
fim FAN_N2558_0 ( .fault(fault), .net(N2558), .FEN(FEN[1363]), .op(N2558_t0) );
fim FAN_N2558_1 ( .fault(fault), .net(N2558), .FEN(FEN[1364]), .op(N2558_t1) );
fim FAN_N2493_0 ( .fault(fault), .net(N2493), .FEN(FEN[1365]), .op(N2493_t0) );
fim FAN_N2493_1 ( .fault(fault), .net(N2493), .FEN(FEN[1366]), .op(N2493_t1) );
fim FAN_N2561_0 ( .fault(fault), .net(N2561), .FEN(FEN[1367]), .op(N2561_t0) );
fim FAN_N2561_1 ( .fault(fault), .net(N2561), .FEN(FEN[1368]), .op(N2561_t1) );
fim FAN_N2498_0 ( .fault(fault), .net(N2498), .FEN(FEN[1369]), .op(N2498_t0) );
fim FAN_N2498_1 ( .fault(fault), .net(N2498), .FEN(FEN[1370]), .op(N2498_t1) );
fim FAN_N2564_0 ( .fault(fault), .net(N2564), .FEN(FEN[1371]), .op(N2564_t0) );
fim FAN_N2564_1 ( .fault(fault), .net(N2564), .FEN(FEN[1372]), .op(N2564_t1) );
fim FAN_N2503_0 ( .fault(fault), .net(N2503), .FEN(FEN[1373]), .op(N2503_t0) );
fim FAN_N2503_1 ( .fault(fault), .net(N2503), .FEN(FEN[1374]), .op(N2503_t1) );
fim FAN_N2567_0 ( .fault(fault), .net(N2567), .FEN(FEN[1375]), .op(N2567_t0) );
fim FAN_N2567_1 ( .fault(fault), .net(N2567), .FEN(FEN[1376]), .op(N2567_t1) );
fim FAN_N2508_0 ( .fault(fault), .net(N2508), .FEN(FEN[1377]), .op(N2508_t0) );
fim FAN_N2508_1 ( .fault(fault), .net(N2508), .FEN(FEN[1378]), .op(N2508_t1) );
fim FAN_N2570_0 ( .fault(fault), .net(N2570), .FEN(FEN[1379]), .op(N2570_t0) );
fim FAN_N2570_1 ( .fault(fault), .net(N2570), .FEN(FEN[1380]), .op(N2570_t1) );
fim FAN_N2513_0 ( .fault(fault), .net(N2513), .FEN(FEN[1381]), .op(N2513_t0) );
fim FAN_N2513_1 ( .fault(fault), .net(N2513), .FEN(FEN[1382]), .op(N2513_t1) );
fim FAN_N2573_0 ( .fault(fault), .net(N2573), .FEN(FEN[1383]), .op(N2573_t0) );
fim FAN_N2573_1 ( .fault(fault), .net(N2573), .FEN(FEN[1384]), .op(N2573_t1) );
fim FAN_N2518_0 ( .fault(fault), .net(N2518), .FEN(FEN[1385]), .op(N2518_t0) );
fim FAN_N2518_1 ( .fault(fault), .net(N2518), .FEN(FEN[1386]), .op(N2518_t1) );
fim FAN_N2576_0 ( .fault(fault), .net(N2576), .FEN(FEN[1387]), .op(N2576_t0) );
fim FAN_N2576_1 ( .fault(fault), .net(N2576), .FEN(FEN[1388]), .op(N2576_t1) );
fim FAN_N2523_0 ( .fault(fault), .net(N2523), .FEN(FEN[1389]), .op(N2523_t0) );
fim FAN_N2523_1 ( .fault(fault), .net(N2523), .FEN(FEN[1390]), .op(N2523_t1) );
fim FAN_N2579_0 ( .fault(fault), .net(N2579), .FEN(FEN[1391]), .op(N2579_t0) );
fim FAN_N2579_1 ( .fault(fault), .net(N2579), .FEN(FEN[1392]), .op(N2579_t1) );
fim FAN_N2528_0 ( .fault(fault), .net(N2528), .FEN(FEN[1393]), .op(N2528_t0) );
fim FAN_N2528_1 ( .fault(fault), .net(N2528), .FEN(FEN[1394]), .op(N2528_t1) );
fim FAN_N2582_0 ( .fault(fault), .net(N2582), .FEN(FEN[1395]), .op(N2582_t0) );
fim FAN_N2582_1 ( .fault(fault), .net(N2582), .FEN(FEN[1396]), .op(N2582_t1) );
fim FAN_N2582_2 ( .fault(fault), .net(N2582), .FEN(FEN[1397]), .op(N2582_t2) );
fim FAN_N2588_0 ( .fault(fault), .net(N2588), .FEN(FEN[1398]), .op(N2588_t0) );
fim FAN_N2588_1 ( .fault(fault), .net(N2588), .FEN(FEN[1399]), .op(N2588_t1) );
fim FAN_N1182_0 ( .fault(fault), .net(N1182), .FEN(FEN[1400]), .op(N1182_t0) );
fim FAN_N1182_1 ( .fault(fault), .net(N1182), .FEN(FEN[1401]), .op(N1182_t1) );
fim FAN_N2591_0 ( .fault(fault), .net(N2591), .FEN(FEN[1402]), .op(N2591_t0) );
fim FAN_N2591_1 ( .fault(fault), .net(N2591), .FEN(FEN[1403]), .op(N2591_t1) );
fim FAN_N2591_2 ( .fault(fault), .net(N2591), .FEN(FEN[1404]), .op(N2591_t2) );
fim FAN_N2595_0 ( .fault(fault), .net(N2595), .FEN(FEN[1405]), .op(N2595_t0) );
fim FAN_N2595_1 ( .fault(fault), .net(N2595), .FEN(FEN[1406]), .op(N2595_t1) );
fim FAN_N2595_2 ( .fault(fault), .net(N2595), .FEN(FEN[1407]), .op(N2595_t2) );
fim FAN_N2599_0 ( .fault(fault), .net(N2599), .FEN(FEN[1408]), .op(N2599_t0) );
fim FAN_N2599_1 ( .fault(fault), .net(N2599), .FEN(FEN[1409]), .op(N2599_t1) );
fim FAN_N2599_2 ( .fault(fault), .net(N2599), .FEN(FEN[1410]), .op(N2599_t2) );
fim FAN_N2603_0 ( .fault(fault), .net(N2603), .FEN(FEN[1411]), .op(N2603_t0) );
fim FAN_N2603_1 ( .fault(fault), .net(N2603), .FEN(FEN[1412]), .op(N2603_t1) );
fim FAN_N2603_2 ( .fault(fault), .net(N2603), .FEN(FEN[1413]), .op(N2603_t2) );
fim FAN_N2607_0 ( .fault(fault), .net(N2607), .FEN(FEN[1414]), .op(N2607_t0) );
fim FAN_N2607_1 ( .fault(fault), .net(N2607), .FEN(FEN[1415]), .op(N2607_t1) );
fim FAN_N2607_2 ( .fault(fault), .net(N2607), .FEN(FEN[1416]), .op(N2607_t2) );
fim FAN_N2611_0 ( .fault(fault), .net(N2611), .FEN(FEN[1417]), .op(N2611_t0) );
fim FAN_N2611_1 ( .fault(fault), .net(N2611), .FEN(FEN[1418]), .op(N2611_t1) );
fim FAN_N2611_2 ( .fault(fault), .net(N2611), .FEN(FEN[1419]), .op(N2611_t2) );
fim FAN_N2615_0 ( .fault(fault), .net(N2615), .FEN(FEN[1420]), .op(N2615_t0) );
fim FAN_N2615_1 ( .fault(fault), .net(N2615), .FEN(FEN[1421]), .op(N2615_t1) );
fim FAN_N2615_2 ( .fault(fault), .net(N2615), .FEN(FEN[1422]), .op(N2615_t2) );
fim FAN_N2619_0 ( .fault(fault), .net(N2619), .FEN(FEN[1423]), .op(N2619_t0) );
fim FAN_N2619_1 ( .fault(fault), .net(N2619), .FEN(FEN[1424]), .op(N2619_t1) );
fim FAN_N2619_2 ( .fault(fault), .net(N2619), .FEN(FEN[1425]), .op(N2619_t2) );
fim FAN_N2623_0 ( .fault(fault), .net(N2623), .FEN(FEN[1426]), .op(N2623_t0) );
fim FAN_N2623_1 ( .fault(fault), .net(N2623), .FEN(FEN[1427]), .op(N2623_t1) );
fim FAN_N2623_2 ( .fault(fault), .net(N2623), .FEN(FEN[1428]), .op(N2623_t2) );
fim FAN_N2627_0 ( .fault(fault), .net(N2627), .FEN(FEN[1429]), .op(N2627_t0) );
fim FAN_N2627_1 ( .fault(fault), .net(N2627), .FEN(FEN[1430]), .op(N2627_t1) );
fim FAN_N2627_2 ( .fault(fault), .net(N2627), .FEN(FEN[1431]), .op(N2627_t2) );
fim FAN_N2631_0 ( .fault(fault), .net(N2631), .FEN(FEN[1432]), .op(N2631_t0) );
fim FAN_N2631_1 ( .fault(fault), .net(N2631), .FEN(FEN[1433]), .op(N2631_t1) );
fim FAN_N2631_2 ( .fault(fault), .net(N2631), .FEN(FEN[1434]), .op(N2631_t2) );
fim FAN_N2635_0 ( .fault(fault), .net(N2635), .FEN(FEN[1435]), .op(N2635_t0) );
fim FAN_N2635_1 ( .fault(fault), .net(N2635), .FEN(FEN[1436]), .op(N2635_t1) );
fim FAN_N2635_2 ( .fault(fault), .net(N2635), .FEN(FEN[1437]), .op(N2635_t2) );
fim FAN_N2641_0 ( .fault(fault), .net(N2641), .FEN(FEN[1438]), .op(N2641_t0) );
fim FAN_N2641_1 ( .fault(fault), .net(N2641), .FEN(FEN[1439]), .op(N2641_t1) );
fim FAN_N1134_0 ( .fault(fault), .net(N1134), .FEN(FEN[1440]), .op(N1134_t0) );
fim FAN_N1134_1 ( .fault(fault), .net(N1134), .FEN(FEN[1441]), .op(N1134_t1) );
fim FAN_N2644_0 ( .fault(fault), .net(N2644), .FEN(FEN[1442]), .op(N2644_t0) );
fim FAN_N2644_1 ( .fault(fault), .net(N2644), .FEN(FEN[1443]), .op(N2644_t1) );
fim FAN_N2644_2 ( .fault(fault), .net(N2644), .FEN(FEN[1444]), .op(N2644_t2) );
fim FAN_N1278_0 ( .fault(fault), .net(N1278), .FEN(FEN[1445]), .op(N1278_t0) );
fim FAN_N1278_1 ( .fault(fault), .net(N1278), .FEN(FEN[1446]), .op(N1278_t1) );
fim FAN_N2650_0 ( .fault(fault), .net(N2650), .FEN(FEN[1447]), .op(N2650_t0) );
fim FAN_N2650_1 ( .fault(fault), .net(N2650), .FEN(FEN[1448]), .op(N2650_t1) );
fim FAN_N2675_0 ( .fault(fault), .net(N2675), .FEN(FEN[1449]), .op(N2675_t0) );
fim FAN_N2675_1 ( .fault(fault), .net(N2675), .FEN(FEN[1450]), .op(N2675_t1) );
fim FAN_N1086_0 ( .fault(fault), .net(N1086), .FEN(FEN[1451]), .op(N1086_t0) );
fim FAN_N1086_1 ( .fault(fault), .net(N1086), .FEN(FEN[1452]), .op(N1086_t1) );
fim FAN_N2678_0 ( .fault(fault), .net(N2678), .FEN(FEN[1453]), .op(N2678_t0) );
fim FAN_N2678_1 ( .fault(fault), .net(N2678), .FEN(FEN[1454]), .op(N2678_t1) );
fim FAN_N2678_2 ( .fault(fault), .net(N2678), .FEN(FEN[1455]), .op(N2678_t2) );
fim FAN_N2687_0 ( .fault(fault), .net(N2687), .FEN(FEN[1456]), .op(N2687_t0) );
fim FAN_N2687_1 ( .fault(fault), .net(N2687), .FEN(FEN[1457]), .op(N2687_t1) );
fim FAN_N2684_0 ( .fault(fault), .net(N2684), .FEN(FEN[1458]), .op(N2684_t0) );
fim FAN_N2684_1 ( .fault(fault), .net(N2684), .FEN(FEN[1459]), .op(N2684_t1) );
fim FAN_N2690_0 ( .fault(fault), .net(N2690), .FEN(FEN[1460]), .op(N2690_t0) );
fim FAN_N2690_1 ( .fault(fault), .net(N2690), .FEN(FEN[1461]), .op(N2690_t1) );
fim FAN_N2690_2 ( .fault(fault), .net(N2690), .FEN(FEN[1462]), .op(N2690_t2) );
fim FAN_N2694_0 ( .fault(fault), .net(N2694), .FEN(FEN[1463]), .op(N2694_t0) );
fim FAN_N2694_1 ( .fault(fault), .net(N2694), .FEN(FEN[1464]), .op(N2694_t1) );
fim FAN_N558_0 ( .fault(fault), .net(N558), .FEN(FEN[1465]), .op(N558_t0) );
fim FAN_N558_1 ( .fault(fault), .net(N558), .FEN(FEN[1466]), .op(N558_t1) );
fim FAN_N2697_0 ( .fault(fault), .net(N2697), .FEN(FEN[1467]), .op(N2697_t0) );
fim FAN_N2697_1 ( .fault(fault), .net(N2697), .FEN(FEN[1468]), .op(N2697_t1) );
fim FAN_N606_0 ( .fault(fault), .net(N606), .FEN(FEN[1469]), .op(N606_t0) );
fim FAN_N606_1 ( .fault(fault), .net(N606), .FEN(FEN[1470]), .op(N606_t1) );
fim FAN_N2700_0 ( .fault(fault), .net(N2700), .FEN(FEN[1471]), .op(N2700_t0) );
fim FAN_N2700_1 ( .fault(fault), .net(N2700), .FEN(FEN[1472]), .op(N2700_t1) );
fim FAN_N654_0 ( .fault(fault), .net(N654), .FEN(FEN[1473]), .op(N654_t0) );
fim FAN_N654_1 ( .fault(fault), .net(N654), .FEN(FEN[1474]), .op(N654_t1) );
fim FAN_N2703_0 ( .fault(fault), .net(N2703), .FEN(FEN[1475]), .op(N2703_t0) );
fim FAN_N2703_1 ( .fault(fault), .net(N2703), .FEN(FEN[1476]), .op(N2703_t1) );
fim FAN_N702_0 ( .fault(fault), .net(N702), .FEN(FEN[1477]), .op(N702_t0) );
fim FAN_N702_1 ( .fault(fault), .net(N702), .FEN(FEN[1478]), .op(N702_t1) );
fim FAN_N2706_0 ( .fault(fault), .net(N2706), .FEN(FEN[1479]), .op(N2706_t0) );
fim FAN_N2706_1 ( .fault(fault), .net(N2706), .FEN(FEN[1480]), .op(N2706_t1) );
fim FAN_N750_0 ( .fault(fault), .net(N750), .FEN(FEN[1481]), .op(N750_t0) );
fim FAN_N750_1 ( .fault(fault), .net(N750), .FEN(FEN[1482]), .op(N750_t1) );
fim FAN_N2709_0 ( .fault(fault), .net(N2709), .FEN(FEN[1483]), .op(N2709_t0) );
fim FAN_N2709_1 ( .fault(fault), .net(N2709), .FEN(FEN[1484]), .op(N2709_t1) );
fim FAN_N798_0 ( .fault(fault), .net(N798), .FEN(FEN[1485]), .op(N798_t0) );
fim FAN_N798_1 ( .fault(fault), .net(N798), .FEN(FEN[1486]), .op(N798_t1) );
fim FAN_N2712_0 ( .fault(fault), .net(N2712), .FEN(FEN[1487]), .op(N2712_t0) );
fim FAN_N2712_1 ( .fault(fault), .net(N2712), .FEN(FEN[1488]), .op(N2712_t1) );
fim FAN_N846_0 ( .fault(fault), .net(N846), .FEN(FEN[1489]), .op(N846_t0) );
fim FAN_N846_1 ( .fault(fault), .net(N846), .FEN(FEN[1490]), .op(N846_t1) );
fim FAN_N2715_0 ( .fault(fault), .net(N2715), .FEN(FEN[1491]), .op(N2715_t0) );
fim FAN_N2715_1 ( .fault(fault), .net(N2715), .FEN(FEN[1492]), .op(N2715_t1) );
fim FAN_N894_0 ( .fault(fault), .net(N894), .FEN(FEN[1493]), .op(N894_t0) );
fim FAN_N894_1 ( .fault(fault), .net(N894), .FEN(FEN[1494]), .op(N894_t1) );
fim FAN_N2718_0 ( .fault(fault), .net(N2718), .FEN(FEN[1495]), .op(N2718_t0) );
fim FAN_N2718_1 ( .fault(fault), .net(N2718), .FEN(FEN[1496]), .op(N2718_t1) );
fim FAN_N942_0 ( .fault(fault), .net(N942), .FEN(FEN[1497]), .op(N942_t0) );
fim FAN_N942_1 ( .fault(fault), .net(N942), .FEN(FEN[1498]), .op(N942_t1) );
fim FAN_N2721_0 ( .fault(fault), .net(N2721), .FEN(FEN[1499]), .op(N2721_t0) );
fim FAN_N2721_1 ( .fault(fault), .net(N2721), .FEN(FEN[1500]), .op(N2721_t1) );
fim FAN_N990_0 ( .fault(fault), .net(N990), .FEN(FEN[1501]), .op(N990_t0) );
fim FAN_N990_1 ( .fault(fault), .net(N990), .FEN(FEN[1502]), .op(N990_t1) );
fim FAN_N2724_0 ( .fault(fault), .net(N2724), .FEN(FEN[1503]), .op(N2724_t0) );
fim FAN_N2724_1 ( .fault(fault), .net(N2724), .FEN(FEN[1504]), .op(N2724_t1) );
fim FAN_N1038_0 ( .fault(fault), .net(N1038), .FEN(FEN[1505]), .op(N1038_t0) );
fim FAN_N1038_1 ( .fault(fault), .net(N1038), .FEN(FEN[1506]), .op(N1038_t1) );
fim FAN_N2727_0 ( .fault(fault), .net(N2727), .FEN(FEN[1507]), .op(N2727_t0) );
fim FAN_N2727_1 ( .fault(fault), .net(N2727), .FEN(FEN[1508]), .op(N2727_t1) );
fim FAN_N2727_2 ( .fault(fault), .net(N2727), .FEN(FEN[1509]), .op(N2727_t2) );
fim FAN_N2736_0 ( .fault(fault), .net(N2736), .FEN(FEN[1510]), .op(N2736_t0) );
fim FAN_N2736_1 ( .fault(fault), .net(N2736), .FEN(FEN[1511]), .op(N2736_t1) );
fim FAN_N2733_0 ( .fault(fault), .net(N2733), .FEN(FEN[1512]), .op(N2733_t0) );
fim FAN_N2733_1 ( .fault(fault), .net(N2733), .FEN(FEN[1513]), .op(N2733_t1) );
fim FAN_N2739_0 ( .fault(fault), .net(N2739), .FEN(FEN[1514]), .op(N2739_t0) );
fim FAN_N2739_1 ( .fault(fault), .net(N2739), .FEN(FEN[1515]), .op(N2739_t1) );
fim FAN_N2739_2 ( .fault(fault), .net(N2739), .FEN(FEN[1516]), .op(N2739_t2) );
fim FAN_N2745_0 ( .fault(fault), .net(N2745), .FEN(FEN[1517]), .op(N2745_t0) );
fim FAN_N2745_1 ( .fault(fault), .net(N2745), .FEN(FEN[1518]), .op(N2745_t1) );
fim FAN_N2745_2 ( .fault(fault), .net(N2745), .FEN(FEN[1519]), .op(N2745_t2) );
fim FAN_N2749_0 ( .fault(fault), .net(N2749), .FEN(FEN[1520]), .op(N2749_t0) );
fim FAN_N2749_1 ( .fault(fault), .net(N2749), .FEN(FEN[1521]), .op(N2749_t1) );
fim FAN_N2749_2 ( .fault(fault), .net(N2749), .FEN(FEN[1522]), .op(N2749_t2) );
fim FAN_N2753_0 ( .fault(fault), .net(N2753), .FEN(FEN[1523]), .op(N2753_t0) );
fim FAN_N2753_1 ( .fault(fault), .net(N2753), .FEN(FEN[1524]), .op(N2753_t1) );
fim FAN_N2753_2 ( .fault(fault), .net(N2753), .FEN(FEN[1525]), .op(N2753_t2) );
fim FAN_N2757_0 ( .fault(fault), .net(N2757), .FEN(FEN[1526]), .op(N2757_t0) );
fim FAN_N2757_1 ( .fault(fault), .net(N2757), .FEN(FEN[1527]), .op(N2757_t1) );
fim FAN_N2757_2 ( .fault(fault), .net(N2757), .FEN(FEN[1528]), .op(N2757_t2) );
fim FAN_N2761_0 ( .fault(fault), .net(N2761), .FEN(FEN[1529]), .op(N2761_t0) );
fim FAN_N2761_1 ( .fault(fault), .net(N2761), .FEN(FEN[1530]), .op(N2761_t1) );
fim FAN_N2761_2 ( .fault(fault), .net(N2761), .FEN(FEN[1531]), .op(N2761_t2) );
fim FAN_N2765_0 ( .fault(fault), .net(N2765), .FEN(FEN[1532]), .op(N2765_t0) );
fim FAN_N2765_1 ( .fault(fault), .net(N2765), .FEN(FEN[1533]), .op(N2765_t1) );
fim FAN_N2765_2 ( .fault(fault), .net(N2765), .FEN(FEN[1534]), .op(N2765_t2) );
fim FAN_N2769_0 ( .fault(fault), .net(N2769), .FEN(FEN[1535]), .op(N2769_t0) );
fim FAN_N2769_1 ( .fault(fault), .net(N2769), .FEN(FEN[1536]), .op(N2769_t1) );
fim FAN_N2769_2 ( .fault(fault), .net(N2769), .FEN(FEN[1537]), .op(N2769_t2) );
fim FAN_N2773_0 ( .fault(fault), .net(N2773), .FEN(FEN[1538]), .op(N2773_t0) );
fim FAN_N2773_1 ( .fault(fault), .net(N2773), .FEN(FEN[1539]), .op(N2773_t1) );
fim FAN_N2773_2 ( .fault(fault), .net(N2773), .FEN(FEN[1540]), .op(N2773_t2) );
fim FAN_N2777_0 ( .fault(fault), .net(N2777), .FEN(FEN[1541]), .op(N2777_t0) );
fim FAN_N2777_1 ( .fault(fault), .net(N2777), .FEN(FEN[1542]), .op(N2777_t1) );
fim FAN_N2777_2 ( .fault(fault), .net(N2777), .FEN(FEN[1543]), .op(N2777_t2) );
fim FAN_N2781_0 ( .fault(fault), .net(N2781), .FEN(FEN[1544]), .op(N2781_t0) );
fim FAN_N2781_1 ( .fault(fault), .net(N2781), .FEN(FEN[1545]), .op(N2781_t1) );
fim FAN_N2781_2 ( .fault(fault), .net(N2781), .FEN(FEN[1546]), .op(N2781_t2) );
fim FAN_N2785_0 ( .fault(fault), .net(N2785), .FEN(FEN[1547]), .op(N2785_t0) );
fim FAN_N2785_1 ( .fault(fault), .net(N2785), .FEN(FEN[1548]), .op(N2785_t1) );
fim FAN_N2785_2 ( .fault(fault), .net(N2785), .FEN(FEN[1549]), .op(N2785_t2) );
fim FAN_N2794_0 ( .fault(fault), .net(N2794), .FEN(FEN[1550]), .op(N2794_t0) );
fim FAN_N2794_1 ( .fault(fault), .net(N2794), .FEN(FEN[1551]), .op(N2794_t1) );
fim FAN_N2791_0 ( .fault(fault), .net(N2791), .FEN(FEN[1552]), .op(N2791_t0) );
fim FAN_N2791_1 ( .fault(fault), .net(N2791), .FEN(FEN[1553]), .op(N2791_t1) );
fim FAN_N2797_0 ( .fault(fault), .net(N2797), .FEN(FEN[1554]), .op(N2797_t0) );
fim FAN_N2797_1 ( .fault(fault), .net(N2797), .FEN(FEN[1555]), .op(N2797_t1) );
fim FAN_N2797_2 ( .fault(fault), .net(N2797), .FEN(FEN[1556]), .op(N2797_t2) );
fim FAN_N2803_0 ( .fault(fault), .net(N2803), .FEN(FEN[1557]), .op(N2803_t0) );
fim FAN_N2803_1 ( .fault(fault), .net(N2803), .FEN(FEN[1558]), .op(N2803_t1) );
fim FAN_N1233_0 ( .fault(fault), .net(N1233), .FEN(FEN[1559]), .op(N1233_t0) );
fim FAN_N1233_1 ( .fault(fault), .net(N1233), .FEN(FEN[1560]), .op(N1233_t1) );
fim FAN_N2861_0 ( .fault(fault), .net(N2861), .FEN(FEN[1561]), .op(N2861_t0) );
fim FAN_N2861_1 ( .fault(fault), .net(N2861), .FEN(FEN[1562]), .op(N2861_t1) );
fim FAN_N2858_0 ( .fault(fault), .net(N2858), .FEN(FEN[1563]), .op(N2858_t0) );
fim FAN_N2858_1 ( .fault(fault), .net(N2858), .FEN(FEN[1564]), .op(N2858_t1) );
fim FAN_N2864_0 ( .fault(fault), .net(N2864), .FEN(FEN[1565]), .op(N2864_t0) );
fim FAN_N2864_1 ( .fault(fault), .net(N2864), .FEN(FEN[1566]), .op(N2864_t1) );
fim FAN_N2864_2 ( .fault(fault), .net(N2864), .FEN(FEN[1567]), .op(N2864_t2) );
fim FAN_N2870_0 ( .fault(fault), .net(N2870), .FEN(FEN[1568]), .op(N2870_t0) );
fim FAN_N2870_1 ( .fault(fault), .net(N2870), .FEN(FEN[1569]), .op(N2870_t1) );
fim FAN_N1185_0 ( .fault(fault), .net(N1185), .FEN(FEN[1570]), .op(N1185_t0) );
fim FAN_N1185_1 ( .fault(fault), .net(N1185), .FEN(FEN[1571]), .op(N1185_t1) );
fim FAN_N2873_0 ( .fault(fault), .net(N2873), .FEN(FEN[1572]), .op(N2873_t0) );
fim FAN_N2873_1 ( .fault(fault), .net(N2873), .FEN(FEN[1573]), .op(N2873_t1) );
fim FAN_N2873_2 ( .fault(fault), .net(N2873), .FEN(FEN[1574]), .op(N2873_t2) );
fim FAN_N2878_0 ( .fault(fault), .net(N2878), .FEN(FEN[1575]), .op(N2878_t0) );
fim FAN_N2878_1 ( .fault(fault), .net(N2878), .FEN(FEN[1576]), .op(N2878_t1) );
fim FAN_N2808_0 ( .fault(fault), .net(N2808), .FEN(FEN[1577]), .op(N2808_t0) );
fim FAN_N2808_1 ( .fault(fault), .net(N2808), .FEN(FEN[1578]), .op(N2808_t1) );
fim FAN_N2881_0 ( .fault(fault), .net(N2881), .FEN(FEN[1579]), .op(N2881_t0) );
fim FAN_N2881_1 ( .fault(fault), .net(N2881), .FEN(FEN[1580]), .op(N2881_t1) );
fim FAN_N2813_0 ( .fault(fault), .net(N2813), .FEN(FEN[1581]), .op(N2813_t0) );
fim FAN_N2813_1 ( .fault(fault), .net(N2813), .FEN(FEN[1582]), .op(N2813_t1) );
fim FAN_N2884_0 ( .fault(fault), .net(N2884), .FEN(FEN[1583]), .op(N2884_t0) );
fim FAN_N2884_1 ( .fault(fault), .net(N2884), .FEN(FEN[1584]), .op(N2884_t1) );
fim FAN_N2818_0 ( .fault(fault), .net(N2818), .FEN(FEN[1585]), .op(N2818_t0) );
fim FAN_N2818_1 ( .fault(fault), .net(N2818), .FEN(FEN[1586]), .op(N2818_t1) );
fim FAN_N2887_0 ( .fault(fault), .net(N2887), .FEN(FEN[1587]), .op(N2887_t0) );
fim FAN_N2887_1 ( .fault(fault), .net(N2887), .FEN(FEN[1588]), .op(N2887_t1) );
fim FAN_N2823_0 ( .fault(fault), .net(N2823), .FEN(FEN[1589]), .op(N2823_t0) );
fim FAN_N2823_1 ( .fault(fault), .net(N2823), .FEN(FEN[1590]), .op(N2823_t1) );
fim FAN_N2890_0 ( .fault(fault), .net(N2890), .FEN(FEN[1591]), .op(N2890_t0) );
fim FAN_N2890_1 ( .fault(fault), .net(N2890), .FEN(FEN[1592]), .op(N2890_t1) );
fim FAN_N2828_0 ( .fault(fault), .net(N2828), .FEN(FEN[1593]), .op(N2828_t0) );
fim FAN_N2828_1 ( .fault(fault), .net(N2828), .FEN(FEN[1594]), .op(N2828_t1) );
fim FAN_N2893_0 ( .fault(fault), .net(N2893), .FEN(FEN[1595]), .op(N2893_t0) );
fim FAN_N2893_1 ( .fault(fault), .net(N2893), .FEN(FEN[1596]), .op(N2893_t1) );
fim FAN_N2833_0 ( .fault(fault), .net(N2833), .FEN(FEN[1597]), .op(N2833_t0) );
fim FAN_N2833_1 ( .fault(fault), .net(N2833), .FEN(FEN[1598]), .op(N2833_t1) );
fim FAN_N2896_0 ( .fault(fault), .net(N2896), .FEN(FEN[1599]), .op(N2896_t0) );
fim FAN_N2896_1 ( .fault(fault), .net(N2896), .FEN(FEN[1600]), .op(N2896_t1) );
fim FAN_N2838_0 ( .fault(fault), .net(N2838), .FEN(FEN[1601]), .op(N2838_t0) );
fim FAN_N2838_1 ( .fault(fault), .net(N2838), .FEN(FEN[1602]), .op(N2838_t1) );
fim FAN_N2899_0 ( .fault(fault), .net(N2899), .FEN(FEN[1603]), .op(N2899_t0) );
fim FAN_N2899_1 ( .fault(fault), .net(N2899), .FEN(FEN[1604]), .op(N2899_t1) );
fim FAN_N2843_0 ( .fault(fault), .net(N2843), .FEN(FEN[1605]), .op(N2843_t0) );
fim FAN_N2843_1 ( .fault(fault), .net(N2843), .FEN(FEN[1606]), .op(N2843_t1) );
fim FAN_N2902_0 ( .fault(fault), .net(N2902), .FEN(FEN[1607]), .op(N2902_t0) );
fim FAN_N2902_1 ( .fault(fault), .net(N2902), .FEN(FEN[1608]), .op(N2902_t1) );
fim FAN_N2848_0 ( .fault(fault), .net(N2848), .FEN(FEN[1609]), .op(N2848_t0) );
fim FAN_N2848_1 ( .fault(fault), .net(N2848), .FEN(FEN[1610]), .op(N2848_t1) );
fim FAN_N2905_0 ( .fault(fault), .net(N2905), .FEN(FEN[1611]), .op(N2905_t0) );
fim FAN_N2905_1 ( .fault(fault), .net(N2905), .FEN(FEN[1612]), .op(N2905_t1) );
fim FAN_N2853_0 ( .fault(fault), .net(N2853), .FEN(FEN[1613]), .op(N2853_t0) );
fim FAN_N2853_1 ( .fault(fault), .net(N2853), .FEN(FEN[1614]), .op(N2853_t1) );
fim FAN_N2908_0 ( .fault(fault), .net(N2908), .FEN(FEN[1615]), .op(N2908_t0) );
fim FAN_N2908_1 ( .fault(fault), .net(N2908), .FEN(FEN[1616]), .op(N2908_t1) );
fim FAN_N2908_2 ( .fault(fault), .net(N2908), .FEN(FEN[1617]), .op(N2908_t2) );
fim FAN_N2914_0 ( .fault(fault), .net(N2914), .FEN(FEN[1618]), .op(N2914_t0) );
fim FAN_N2914_1 ( .fault(fault), .net(N2914), .FEN(FEN[1619]), .op(N2914_t1) );
fim FAN_N1137_0 ( .fault(fault), .net(N1137), .FEN(FEN[1620]), .op(N1137_t0) );
fim FAN_N1137_1 ( .fault(fault), .net(N1137), .FEN(FEN[1621]), .op(N1137_t1) );
fim FAN_N2917_0 ( .fault(fault), .net(N2917), .FEN(FEN[1622]), .op(N2917_t0) );
fim FAN_N2917_1 ( .fault(fault), .net(N2917), .FEN(FEN[1623]), .op(N2917_t1) );
fim FAN_N2917_2 ( .fault(fault), .net(N2917), .FEN(FEN[1624]), .op(N2917_t2) );
fim FAN_N1281_0 ( .fault(fault), .net(N1281), .FEN(FEN[1625]), .op(N1281_t0) );
fim FAN_N1281_1 ( .fault(fault), .net(N1281), .FEN(FEN[1626]), .op(N1281_t1) );
fim FAN_N2923_0 ( .fault(fault), .net(N2923), .FEN(FEN[1627]), .op(N2923_t0) );
fim FAN_N2923_1 ( .fault(fault), .net(N2923), .FEN(FEN[1628]), .op(N2923_t1) );
fim FAN_N2926_0 ( .fault(fault), .net(N2926), .FEN(FEN[1629]), .op(N2926_t0) );
fim FAN_N2926_1 ( .fault(fault), .net(N2926), .FEN(FEN[1630]), .op(N2926_t1) );
fim FAN_N2926_2 ( .fault(fault), .net(N2926), .FEN(FEN[1631]), .op(N2926_t2) );
fim FAN_N2930_0 ( .fault(fault), .net(N2930), .FEN(FEN[1632]), .op(N2930_t0) );
fim FAN_N2930_1 ( .fault(fault), .net(N2930), .FEN(FEN[1633]), .op(N2930_t1) );
fim FAN_N2930_2 ( .fault(fault), .net(N2930), .FEN(FEN[1634]), .op(N2930_t2) );
fim FAN_N2934_0 ( .fault(fault), .net(N2934), .FEN(FEN[1635]), .op(N2934_t0) );
fim FAN_N2934_1 ( .fault(fault), .net(N2934), .FEN(FEN[1636]), .op(N2934_t1) );
fim FAN_N2934_2 ( .fault(fault), .net(N2934), .FEN(FEN[1637]), .op(N2934_t2) );
fim FAN_N2938_0 ( .fault(fault), .net(N2938), .FEN(FEN[1638]), .op(N2938_t0) );
fim FAN_N2938_1 ( .fault(fault), .net(N2938), .FEN(FEN[1639]), .op(N2938_t1) );
fim FAN_N2938_2 ( .fault(fault), .net(N2938), .FEN(FEN[1640]), .op(N2938_t2) );
fim FAN_N2942_0 ( .fault(fault), .net(N2942), .FEN(FEN[1641]), .op(N2942_t0) );
fim FAN_N2942_1 ( .fault(fault), .net(N2942), .FEN(FEN[1642]), .op(N2942_t1) );
fim FAN_N2942_2 ( .fault(fault), .net(N2942), .FEN(FEN[1643]), .op(N2942_t2) );
fim FAN_N2946_0 ( .fault(fault), .net(N2946), .FEN(FEN[1644]), .op(N2946_t0) );
fim FAN_N2946_1 ( .fault(fault), .net(N2946), .FEN(FEN[1645]), .op(N2946_t1) );
fim FAN_N2946_2 ( .fault(fault), .net(N2946), .FEN(FEN[1646]), .op(N2946_t2) );
fim FAN_N2950_0 ( .fault(fault), .net(N2950), .FEN(FEN[1647]), .op(N2950_t0) );
fim FAN_N2950_1 ( .fault(fault), .net(N2950), .FEN(FEN[1648]), .op(N2950_t1) );
fim FAN_N2950_2 ( .fault(fault), .net(N2950), .FEN(FEN[1649]), .op(N2950_t2) );
fim FAN_N2954_0 ( .fault(fault), .net(N2954), .FEN(FEN[1650]), .op(N2954_t0) );
fim FAN_N2954_1 ( .fault(fault), .net(N2954), .FEN(FEN[1651]), .op(N2954_t1) );
fim FAN_N2954_2 ( .fault(fault), .net(N2954), .FEN(FEN[1652]), .op(N2954_t2) );
fim FAN_N2958_0 ( .fault(fault), .net(N2958), .FEN(FEN[1653]), .op(N2958_t0) );
fim FAN_N2958_1 ( .fault(fault), .net(N2958), .FEN(FEN[1654]), .op(N2958_t1) );
fim FAN_N2958_2 ( .fault(fault), .net(N2958), .FEN(FEN[1655]), .op(N2958_t2) );
fim FAN_N2962_0 ( .fault(fault), .net(N2962), .FEN(FEN[1656]), .op(N2962_t0) );
fim FAN_N2962_1 ( .fault(fault), .net(N2962), .FEN(FEN[1657]), .op(N2962_t1) );
fim FAN_N2962_2 ( .fault(fault), .net(N2962), .FEN(FEN[1658]), .op(N2962_t2) );
fim FAN_N2968_0 ( .fault(fault), .net(N2968), .FEN(FEN[1659]), .op(N2968_t0) );
fim FAN_N2968_1 ( .fault(fault), .net(N2968), .FEN(FEN[1660]), .op(N2968_t1) );
fim FAN_N1089_0 ( .fault(fault), .net(N1089), .FEN(FEN[1661]), .op(N1089_t0) );
fim FAN_N1089_1 ( .fault(fault), .net(N1089), .FEN(FEN[1662]), .op(N1089_t1) );
fim FAN_N2971_0 ( .fault(fault), .net(N2971), .FEN(FEN[1663]), .op(N2971_t0) );
fim FAN_N2971_1 ( .fault(fault), .net(N2971), .FEN(FEN[1664]), .op(N2971_t1) );
fim FAN_N2971_2 ( .fault(fault), .net(N2971), .FEN(FEN[1665]), .op(N2971_t2) );
fim FAN_N2980_0 ( .fault(fault), .net(N2980), .FEN(FEN[1666]), .op(N2980_t0) );
fim FAN_N2980_1 ( .fault(fault), .net(N2980), .FEN(FEN[1667]), .op(N2980_t1) );
fim FAN_N2977_0 ( .fault(fault), .net(N2977), .FEN(FEN[1668]), .op(N2977_t0) );
fim FAN_N2977_1 ( .fault(fault), .net(N2977), .FEN(FEN[1669]), .op(N2977_t1) );
fim FAN_N2983_0 ( .fault(fault), .net(N2983), .FEN(FEN[1670]), .op(N2983_t0) );
fim FAN_N2983_1 ( .fault(fault), .net(N2983), .FEN(FEN[1671]), .op(N2983_t1) );
fim FAN_N2983_2 ( .fault(fault), .net(N2983), .FEN(FEN[1672]), .op(N2983_t2) );
fim FAN_N3007_0 ( .fault(fault), .net(N3007), .FEN(FEN[1673]), .op(N3007_t0) );
fim FAN_N3007_1 ( .fault(fault), .net(N3007), .FEN(FEN[1674]), .op(N3007_t1) );
fim FAN_N1041_0 ( .fault(fault), .net(N1041), .FEN(FEN[1675]), .op(N1041_t0) );
fim FAN_N1041_1 ( .fault(fault), .net(N1041), .FEN(FEN[1676]), .op(N1041_t1) );
fim FAN_N3010_0 ( .fault(fault), .net(N3010), .FEN(FEN[1677]), .op(N3010_t0) );
fim FAN_N3010_1 ( .fault(fault), .net(N3010), .FEN(FEN[1678]), .op(N3010_t1) );
fim FAN_N3010_2 ( .fault(fault), .net(N3010), .FEN(FEN[1679]), .op(N3010_t2) );
fim FAN_N3019_0 ( .fault(fault), .net(N3019), .FEN(FEN[1680]), .op(N3019_t0) );
fim FAN_N3019_1 ( .fault(fault), .net(N3019), .FEN(FEN[1681]), .op(N3019_t1) );
fim FAN_N3016_0 ( .fault(fault), .net(N3016), .FEN(FEN[1682]), .op(N3016_t0) );
fim FAN_N3016_1 ( .fault(fault), .net(N3016), .FEN(FEN[1683]), .op(N3016_t1) );
fim FAN_N3022_0 ( .fault(fault), .net(N3022), .FEN(FEN[1684]), .op(N3022_t0) );
fim FAN_N3022_1 ( .fault(fault), .net(N3022), .FEN(FEN[1685]), .op(N3022_t1) );
fim FAN_N3022_2 ( .fault(fault), .net(N3022), .FEN(FEN[1686]), .op(N3022_t2) );
fim FAN_N3028_0 ( .fault(fault), .net(N3028), .FEN(FEN[1687]), .op(N3028_t0) );
fim FAN_N3028_1 ( .fault(fault), .net(N3028), .FEN(FEN[1688]), .op(N3028_t1) );
fim FAN_N561_0 ( .fault(fault), .net(N561), .FEN(FEN[1689]), .op(N561_t0) );
fim FAN_N561_1 ( .fault(fault), .net(N561), .FEN(FEN[1690]), .op(N561_t1) );
fim FAN_N3031_0 ( .fault(fault), .net(N3031), .FEN(FEN[1691]), .op(N3031_t0) );
fim FAN_N3031_1 ( .fault(fault), .net(N3031), .FEN(FEN[1692]), .op(N3031_t1) );
fim FAN_N609_0 ( .fault(fault), .net(N609), .FEN(FEN[1693]), .op(N609_t0) );
fim FAN_N609_1 ( .fault(fault), .net(N609), .FEN(FEN[1694]), .op(N609_t1) );
fim FAN_N3034_0 ( .fault(fault), .net(N3034), .FEN(FEN[1695]), .op(N3034_t0) );
fim FAN_N3034_1 ( .fault(fault), .net(N3034), .FEN(FEN[1696]), .op(N3034_t1) );
fim FAN_N657_0 ( .fault(fault), .net(N657), .FEN(FEN[1697]), .op(N657_t0) );
fim FAN_N657_1 ( .fault(fault), .net(N657), .FEN(FEN[1698]), .op(N657_t1) );
fim FAN_N3037_0 ( .fault(fault), .net(N3037), .FEN(FEN[1699]), .op(N3037_t0) );
fim FAN_N3037_1 ( .fault(fault), .net(N3037), .FEN(FEN[1700]), .op(N3037_t1) );
fim FAN_N705_0 ( .fault(fault), .net(N705), .FEN(FEN[1701]), .op(N705_t0) );
fim FAN_N705_1 ( .fault(fault), .net(N705), .FEN(FEN[1702]), .op(N705_t1) );
fim FAN_N3040_0 ( .fault(fault), .net(N3040), .FEN(FEN[1703]), .op(N3040_t0) );
fim FAN_N3040_1 ( .fault(fault), .net(N3040), .FEN(FEN[1704]), .op(N3040_t1) );
fim FAN_N753_0 ( .fault(fault), .net(N753), .FEN(FEN[1705]), .op(N753_t0) );
fim FAN_N753_1 ( .fault(fault), .net(N753), .FEN(FEN[1706]), .op(N753_t1) );
fim FAN_N3043_0 ( .fault(fault), .net(N3043), .FEN(FEN[1707]), .op(N3043_t0) );
fim FAN_N3043_1 ( .fault(fault), .net(N3043), .FEN(FEN[1708]), .op(N3043_t1) );
fim FAN_N801_0 ( .fault(fault), .net(N801), .FEN(FEN[1709]), .op(N801_t0) );
fim FAN_N801_1 ( .fault(fault), .net(N801), .FEN(FEN[1710]), .op(N801_t1) );
fim FAN_N3046_0 ( .fault(fault), .net(N3046), .FEN(FEN[1711]), .op(N3046_t0) );
fim FAN_N3046_1 ( .fault(fault), .net(N3046), .FEN(FEN[1712]), .op(N3046_t1) );
fim FAN_N849_0 ( .fault(fault), .net(N849), .FEN(FEN[1713]), .op(N849_t0) );
fim FAN_N849_1 ( .fault(fault), .net(N849), .FEN(FEN[1714]), .op(N849_t1) );
fim FAN_N3049_0 ( .fault(fault), .net(N3049), .FEN(FEN[1715]), .op(N3049_t0) );
fim FAN_N3049_1 ( .fault(fault), .net(N3049), .FEN(FEN[1716]), .op(N3049_t1) );
fim FAN_N897_0 ( .fault(fault), .net(N897), .FEN(FEN[1717]), .op(N897_t0) );
fim FAN_N897_1 ( .fault(fault), .net(N897), .FEN(FEN[1718]), .op(N897_t1) );
fim FAN_N3052_0 ( .fault(fault), .net(N3052), .FEN(FEN[1719]), .op(N3052_t0) );
fim FAN_N3052_1 ( .fault(fault), .net(N3052), .FEN(FEN[1720]), .op(N3052_t1) );
fim FAN_N945_0 ( .fault(fault), .net(N945), .FEN(FEN[1721]), .op(N945_t0) );
fim FAN_N945_1 ( .fault(fault), .net(N945), .FEN(FEN[1722]), .op(N945_t1) );
fim FAN_N3055_0 ( .fault(fault), .net(N3055), .FEN(FEN[1723]), .op(N3055_t0) );
fim FAN_N3055_1 ( .fault(fault), .net(N3055), .FEN(FEN[1724]), .op(N3055_t1) );
fim FAN_N993_0 ( .fault(fault), .net(N993), .FEN(FEN[1725]), .op(N993_t0) );
fim FAN_N993_1 ( .fault(fault), .net(N993), .FEN(FEN[1726]), .op(N993_t1) );
fim FAN_N3058_0 ( .fault(fault), .net(N3058), .FEN(FEN[1727]), .op(N3058_t0) );
fim FAN_N3058_1 ( .fault(fault), .net(N3058), .FEN(FEN[1728]), .op(N3058_t1) );
fim FAN_N3058_2 ( .fault(fault), .net(N3058), .FEN(FEN[1729]), .op(N3058_t2) );
fim FAN_N3067_0 ( .fault(fault), .net(N3067), .FEN(FEN[1730]), .op(N3067_t0) );
fim FAN_N3067_1 ( .fault(fault), .net(N3067), .FEN(FEN[1731]), .op(N3067_t1) );
fim FAN_N3064_0 ( .fault(fault), .net(N3064), .FEN(FEN[1732]), .op(N3064_t0) );
fim FAN_N3064_1 ( .fault(fault), .net(N3064), .FEN(FEN[1733]), .op(N3064_t1) );
fim FAN_N3070_0 ( .fault(fault), .net(N3070), .FEN(FEN[1734]), .op(N3070_t0) );
fim FAN_N3070_1 ( .fault(fault), .net(N3070), .FEN(FEN[1735]), .op(N3070_t1) );
fim FAN_N3070_2 ( .fault(fault), .net(N3070), .FEN(FEN[1736]), .op(N3070_t2) );
fim FAN_N3076_0 ( .fault(fault), .net(N3076), .FEN(FEN[1737]), .op(N3076_t0) );
fim FAN_N3076_1 ( .fault(fault), .net(N3076), .FEN(FEN[1738]), .op(N3076_t1) );
fim FAN_N1236_0 ( .fault(fault), .net(N1236), .FEN(FEN[1739]), .op(N1236_t0) );
fim FAN_N1236_1 ( .fault(fault), .net(N1236), .FEN(FEN[1740]), .op(N1236_t1) );
fim FAN_N3079_0 ( .fault(fault), .net(N3079), .FEN(FEN[1741]), .op(N3079_t0) );
fim FAN_N3079_1 ( .fault(fault), .net(N3079), .FEN(FEN[1742]), .op(N3079_t1) );
fim FAN_N3079_2 ( .fault(fault), .net(N3079), .FEN(FEN[1743]), .op(N3079_t2) );
fim FAN_N3083_0 ( .fault(fault), .net(N3083), .FEN(FEN[1744]), .op(N3083_t0) );
fim FAN_N3083_1 ( .fault(fault), .net(N3083), .FEN(FEN[1745]), .op(N3083_t1) );
fim FAN_N3083_2 ( .fault(fault), .net(N3083), .FEN(FEN[1746]), .op(N3083_t2) );
fim FAN_N3087_0 ( .fault(fault), .net(N3087), .FEN(FEN[1747]), .op(N3087_t0) );
fim FAN_N3087_1 ( .fault(fault), .net(N3087), .FEN(FEN[1748]), .op(N3087_t1) );
fim FAN_N3087_2 ( .fault(fault), .net(N3087), .FEN(FEN[1749]), .op(N3087_t2) );
fim FAN_N3091_0 ( .fault(fault), .net(N3091), .FEN(FEN[1750]), .op(N3091_t0) );
fim FAN_N3091_1 ( .fault(fault), .net(N3091), .FEN(FEN[1751]), .op(N3091_t1) );
fim FAN_N3091_2 ( .fault(fault), .net(N3091), .FEN(FEN[1752]), .op(N3091_t2) );
fim FAN_N3095_0 ( .fault(fault), .net(N3095), .FEN(FEN[1753]), .op(N3095_t0) );
fim FAN_N3095_1 ( .fault(fault), .net(N3095), .FEN(FEN[1754]), .op(N3095_t1) );
fim FAN_N3095_2 ( .fault(fault), .net(N3095), .FEN(FEN[1755]), .op(N3095_t2) );
fim FAN_N3099_0 ( .fault(fault), .net(N3099), .FEN(FEN[1756]), .op(N3099_t0) );
fim FAN_N3099_1 ( .fault(fault), .net(N3099), .FEN(FEN[1757]), .op(N3099_t1) );
fim FAN_N3099_2 ( .fault(fault), .net(N3099), .FEN(FEN[1758]), .op(N3099_t2) );
fim FAN_N3103_0 ( .fault(fault), .net(N3103), .FEN(FEN[1759]), .op(N3103_t0) );
fim FAN_N3103_1 ( .fault(fault), .net(N3103), .FEN(FEN[1760]), .op(N3103_t1) );
fim FAN_N3103_2 ( .fault(fault), .net(N3103), .FEN(FEN[1761]), .op(N3103_t2) );
fim FAN_N3107_0 ( .fault(fault), .net(N3107), .FEN(FEN[1762]), .op(N3107_t0) );
fim FAN_N3107_1 ( .fault(fault), .net(N3107), .FEN(FEN[1763]), .op(N3107_t1) );
fim FAN_N3107_2 ( .fault(fault), .net(N3107), .FEN(FEN[1764]), .op(N3107_t2) );
fim FAN_N3111_0 ( .fault(fault), .net(N3111), .FEN(FEN[1765]), .op(N3111_t0) );
fim FAN_N3111_1 ( .fault(fault), .net(N3111), .FEN(FEN[1766]), .op(N3111_t1) );
fim FAN_N3111_2 ( .fault(fault), .net(N3111), .FEN(FEN[1767]), .op(N3111_t2) );
fim FAN_N3115_0 ( .fault(fault), .net(N3115), .FEN(FEN[1768]), .op(N3115_t0) );
fim FAN_N3115_1 ( .fault(fault), .net(N3115), .FEN(FEN[1769]), .op(N3115_t1) );
fim FAN_N3115_2 ( .fault(fault), .net(N3115), .FEN(FEN[1770]), .op(N3115_t2) );
fim FAN_N3124_0 ( .fault(fault), .net(N3124), .FEN(FEN[1771]), .op(N3124_t0) );
fim FAN_N3124_1 ( .fault(fault), .net(N3124), .FEN(FEN[1772]), .op(N3124_t1) );
fim FAN_N3121_0 ( .fault(fault), .net(N3121), .FEN(FEN[1773]), .op(N3121_t0) );
fim FAN_N3121_1 ( .fault(fault), .net(N3121), .FEN(FEN[1774]), .op(N3121_t1) );
fim FAN_N3127_0 ( .fault(fault), .net(N3127), .FEN(FEN[1775]), .op(N3127_t0) );
fim FAN_N3127_1 ( .fault(fault), .net(N3127), .FEN(FEN[1776]), .op(N3127_t1) );
fim FAN_N3127_2 ( .fault(fault), .net(N3127), .FEN(FEN[1777]), .op(N3127_t2) );
fim FAN_N3133_0 ( .fault(fault), .net(N3133), .FEN(FEN[1778]), .op(N3133_t0) );
fim FAN_N3133_1 ( .fault(fault), .net(N3133), .FEN(FEN[1779]), .op(N3133_t1) );
fim FAN_N1188_0 ( .fault(fault), .net(N1188), .FEN(FEN[1780]), .op(N1188_t0) );
fim FAN_N1188_1 ( .fault(fault), .net(N1188), .FEN(FEN[1781]), .op(N1188_t1) );
fim FAN_N3136_0 ( .fault(fault), .net(N3136), .FEN(FEN[1782]), .op(N3136_t0) );
fim FAN_N3136_1 ( .fault(fault), .net(N3136), .FEN(FEN[1783]), .op(N3136_t1) );
fim FAN_N3136_2 ( .fault(fault), .net(N3136), .FEN(FEN[1784]), .op(N3136_t2) );
fim FAN_N3190_0 ( .fault(fault), .net(N3190), .FEN(FEN[1785]), .op(N3190_t0) );
fim FAN_N3190_1 ( .fault(fault), .net(N3190), .FEN(FEN[1786]), .op(N3190_t1) );
fim FAN_N3187_0 ( .fault(fault), .net(N3187), .FEN(FEN[1787]), .op(N3187_t0) );
fim FAN_N3187_1 ( .fault(fault), .net(N3187), .FEN(FEN[1788]), .op(N3187_t1) );
fim FAN_N3193_0 ( .fault(fault), .net(N3193), .FEN(FEN[1789]), .op(N3193_t0) );
fim FAN_N3193_1 ( .fault(fault), .net(N3193), .FEN(FEN[1790]), .op(N3193_t1) );
fim FAN_N3193_2 ( .fault(fault), .net(N3193), .FEN(FEN[1791]), .op(N3193_t2) );
fim FAN_N3199_0 ( .fault(fault), .net(N3199), .FEN(FEN[1792]), .op(N3199_t0) );
fim FAN_N3199_1 ( .fault(fault), .net(N3199), .FEN(FEN[1793]), .op(N3199_t1) );
fim FAN_N1140_0 ( .fault(fault), .net(N1140), .FEN(FEN[1794]), .op(N1140_t0) );
fim FAN_N1140_1 ( .fault(fault), .net(N1140), .FEN(FEN[1795]), .op(N1140_t1) );
fim FAN_N3202_0 ( .fault(fault), .net(N3202), .FEN(FEN[1796]), .op(N3202_t0) );
fim FAN_N3202_1 ( .fault(fault), .net(N3202), .FEN(FEN[1797]), .op(N3202_t1) );
fim FAN_N3202_2 ( .fault(fault), .net(N3202), .FEN(FEN[1798]), .op(N3202_t2) );
fim FAN_N1284_0 ( .fault(fault), .net(N1284), .FEN(FEN[1799]), .op(N1284_t0) );
fim FAN_N1284_1 ( .fault(fault), .net(N1284), .FEN(FEN[1800]), .op(N1284_t1) );
fim FAN_N3208_0 ( .fault(fault), .net(N3208), .FEN(FEN[1801]), .op(N3208_t0) );
fim FAN_N3208_1 ( .fault(fault), .net(N3208), .FEN(FEN[1802]), .op(N3208_t1) );
fim FAN_N3212_0 ( .fault(fault), .net(N3212), .FEN(FEN[1803]), .op(N3212_t0) );
fim FAN_N3212_1 ( .fault(fault), .net(N3212), .FEN(FEN[1804]), .op(N3212_t1) );
fim FAN_N3142_0 ( .fault(fault), .net(N3142), .FEN(FEN[1805]), .op(N3142_t0) );
fim FAN_N3142_1 ( .fault(fault), .net(N3142), .FEN(FEN[1806]), .op(N3142_t1) );
fim FAN_N3215_0 ( .fault(fault), .net(N3215), .FEN(FEN[1807]), .op(N3215_t0) );
fim FAN_N3215_1 ( .fault(fault), .net(N3215), .FEN(FEN[1808]), .op(N3215_t1) );
fim FAN_N3147_0 ( .fault(fault), .net(N3147), .FEN(FEN[1809]), .op(N3147_t0) );
fim FAN_N3147_1 ( .fault(fault), .net(N3147), .FEN(FEN[1810]), .op(N3147_t1) );
fim FAN_N3218_0 ( .fault(fault), .net(N3218), .FEN(FEN[1811]), .op(N3218_t0) );
fim FAN_N3218_1 ( .fault(fault), .net(N3218), .FEN(FEN[1812]), .op(N3218_t1) );
fim FAN_N3152_0 ( .fault(fault), .net(N3152), .FEN(FEN[1813]), .op(N3152_t0) );
fim FAN_N3152_1 ( .fault(fault), .net(N3152), .FEN(FEN[1814]), .op(N3152_t1) );
fim FAN_N3221_0 ( .fault(fault), .net(N3221), .FEN(FEN[1815]), .op(N3221_t0) );
fim FAN_N3221_1 ( .fault(fault), .net(N3221), .FEN(FEN[1816]), .op(N3221_t1) );
fim FAN_N3157_0 ( .fault(fault), .net(N3157), .FEN(FEN[1817]), .op(N3157_t0) );
fim FAN_N3157_1 ( .fault(fault), .net(N3157), .FEN(FEN[1818]), .op(N3157_t1) );
fim FAN_N3224_0 ( .fault(fault), .net(N3224), .FEN(FEN[1819]), .op(N3224_t0) );
fim FAN_N3224_1 ( .fault(fault), .net(N3224), .FEN(FEN[1820]), .op(N3224_t1) );
fim FAN_N3162_0 ( .fault(fault), .net(N3162), .FEN(FEN[1821]), .op(N3162_t0) );
fim FAN_N3162_1 ( .fault(fault), .net(N3162), .FEN(FEN[1822]), .op(N3162_t1) );
fim FAN_N3227_0 ( .fault(fault), .net(N3227), .FEN(FEN[1823]), .op(N3227_t0) );
fim FAN_N3227_1 ( .fault(fault), .net(N3227), .FEN(FEN[1824]), .op(N3227_t1) );
fim FAN_N3167_0 ( .fault(fault), .net(N3167), .FEN(FEN[1825]), .op(N3167_t0) );
fim FAN_N3167_1 ( .fault(fault), .net(N3167), .FEN(FEN[1826]), .op(N3167_t1) );
fim FAN_N3230_0 ( .fault(fault), .net(N3230), .FEN(FEN[1827]), .op(N3230_t0) );
fim FAN_N3230_1 ( .fault(fault), .net(N3230), .FEN(FEN[1828]), .op(N3230_t1) );
fim FAN_N3172_0 ( .fault(fault), .net(N3172), .FEN(FEN[1829]), .op(N3172_t0) );
fim FAN_N3172_1 ( .fault(fault), .net(N3172), .FEN(FEN[1830]), .op(N3172_t1) );
fim FAN_N3233_0 ( .fault(fault), .net(N3233), .FEN(FEN[1831]), .op(N3233_t0) );
fim FAN_N3233_1 ( .fault(fault), .net(N3233), .FEN(FEN[1832]), .op(N3233_t1) );
fim FAN_N3177_0 ( .fault(fault), .net(N3177), .FEN(FEN[1833]), .op(N3177_t0) );
fim FAN_N3177_1 ( .fault(fault), .net(N3177), .FEN(FEN[1834]), .op(N3177_t1) );
fim FAN_N3236_0 ( .fault(fault), .net(N3236), .FEN(FEN[1835]), .op(N3236_t0) );
fim FAN_N3236_1 ( .fault(fault), .net(N3236), .FEN(FEN[1836]), .op(N3236_t1) );
fim FAN_N3182_0 ( .fault(fault), .net(N3182), .FEN(FEN[1837]), .op(N3182_t0) );
fim FAN_N3182_1 ( .fault(fault), .net(N3182), .FEN(FEN[1838]), .op(N3182_t1) );
fim FAN_N3239_0 ( .fault(fault), .net(N3239), .FEN(FEN[1839]), .op(N3239_t0) );
fim FAN_N3239_1 ( .fault(fault), .net(N3239), .FEN(FEN[1840]), .op(N3239_t1) );
fim FAN_N3239_2 ( .fault(fault), .net(N3239), .FEN(FEN[1841]), .op(N3239_t2) );
fim FAN_N3245_0 ( .fault(fault), .net(N3245), .FEN(FEN[1842]), .op(N3245_t0) );
fim FAN_N3245_1 ( .fault(fault), .net(N3245), .FEN(FEN[1843]), .op(N3245_t1) );
fim FAN_N1092_0 ( .fault(fault), .net(N1092), .FEN(FEN[1844]), .op(N1092_t0) );
fim FAN_N1092_1 ( .fault(fault), .net(N1092), .FEN(FEN[1845]), .op(N1092_t1) );
fim FAN_N3248_0 ( .fault(fault), .net(N3248), .FEN(FEN[1846]), .op(N3248_t0) );
fim FAN_N3248_1 ( .fault(fault), .net(N3248), .FEN(FEN[1847]), .op(N3248_t1) );
fim FAN_N3248_2 ( .fault(fault), .net(N3248), .FEN(FEN[1848]), .op(N3248_t2) );
fim FAN_N3257_0 ( .fault(fault), .net(N3257), .FEN(FEN[1849]), .op(N3257_t0) );
fim FAN_N3257_1 ( .fault(fault), .net(N3257), .FEN(FEN[1850]), .op(N3257_t1) );
fim FAN_N3254_0 ( .fault(fault), .net(N3254), .FEN(FEN[1851]), .op(N3254_t0) );
fim FAN_N3254_1 ( .fault(fault), .net(N3254), .FEN(FEN[1852]), .op(N3254_t1) );
fim FAN_N3260_0 ( .fault(fault), .net(N3260), .FEN(FEN[1853]), .op(N3260_t0) );
fim FAN_N3260_1 ( .fault(fault), .net(N3260), .FEN(FEN[1854]), .op(N3260_t1) );
fim FAN_N3260_2 ( .fault(fault), .net(N3260), .FEN(FEN[1855]), .op(N3260_t2) );
fim FAN_N3264_0 ( .fault(fault), .net(N3264), .FEN(FEN[1856]), .op(N3264_t0) );
fim FAN_N3264_1 ( .fault(fault), .net(N3264), .FEN(FEN[1857]), .op(N3264_t1) );
fim FAN_N3264_2 ( .fault(fault), .net(N3264), .FEN(FEN[1858]), .op(N3264_t2) );
fim FAN_N3268_0 ( .fault(fault), .net(N3268), .FEN(FEN[1859]), .op(N3268_t0) );
fim FAN_N3268_1 ( .fault(fault), .net(N3268), .FEN(FEN[1860]), .op(N3268_t1) );
fim FAN_N3268_2 ( .fault(fault), .net(N3268), .FEN(FEN[1861]), .op(N3268_t2) );
fim FAN_N3272_0 ( .fault(fault), .net(N3272), .FEN(FEN[1862]), .op(N3272_t0) );
fim FAN_N3272_1 ( .fault(fault), .net(N3272), .FEN(FEN[1863]), .op(N3272_t1) );
fim FAN_N3272_2 ( .fault(fault), .net(N3272), .FEN(FEN[1864]), .op(N3272_t2) );
fim FAN_N3276_0 ( .fault(fault), .net(N3276), .FEN(FEN[1865]), .op(N3276_t0) );
fim FAN_N3276_1 ( .fault(fault), .net(N3276), .FEN(FEN[1866]), .op(N3276_t1) );
fim FAN_N3276_2 ( .fault(fault), .net(N3276), .FEN(FEN[1867]), .op(N3276_t2) );
fim FAN_N3280_0 ( .fault(fault), .net(N3280), .FEN(FEN[1868]), .op(N3280_t0) );
fim FAN_N3280_1 ( .fault(fault), .net(N3280), .FEN(FEN[1869]), .op(N3280_t1) );
fim FAN_N3280_2 ( .fault(fault), .net(N3280), .FEN(FEN[1870]), .op(N3280_t2) );
fim FAN_N3284_0 ( .fault(fault), .net(N3284), .FEN(FEN[1871]), .op(N3284_t0) );
fim FAN_N3284_1 ( .fault(fault), .net(N3284), .FEN(FEN[1872]), .op(N3284_t1) );
fim FAN_N3284_2 ( .fault(fault), .net(N3284), .FEN(FEN[1873]), .op(N3284_t2) );
fim FAN_N3288_0 ( .fault(fault), .net(N3288), .FEN(FEN[1874]), .op(N3288_t0) );
fim FAN_N3288_1 ( .fault(fault), .net(N3288), .FEN(FEN[1875]), .op(N3288_t1) );
fim FAN_N3288_2 ( .fault(fault), .net(N3288), .FEN(FEN[1876]), .op(N3288_t2) );
fim FAN_N3292_0 ( .fault(fault), .net(N3292), .FEN(FEN[1877]), .op(N3292_t0) );
fim FAN_N3292_1 ( .fault(fault), .net(N3292), .FEN(FEN[1878]), .op(N3292_t1) );
fim FAN_N3292_2 ( .fault(fault), .net(N3292), .FEN(FEN[1879]), .op(N3292_t2) );
fim FAN_N3296_0 ( .fault(fault), .net(N3296), .FEN(FEN[1880]), .op(N3296_t0) );
fim FAN_N3296_1 ( .fault(fault), .net(N3296), .FEN(FEN[1881]), .op(N3296_t1) );
fim FAN_N3296_2 ( .fault(fault), .net(N3296), .FEN(FEN[1882]), .op(N3296_t2) );
fim FAN_N3302_0 ( .fault(fault), .net(N3302), .FEN(FEN[1883]), .op(N3302_t0) );
fim FAN_N3302_1 ( .fault(fault), .net(N3302), .FEN(FEN[1884]), .op(N3302_t1) );
fim FAN_N1044_0 ( .fault(fault), .net(N1044), .FEN(FEN[1885]), .op(N1044_t0) );
fim FAN_N1044_1 ( .fault(fault), .net(N1044), .FEN(FEN[1886]), .op(N1044_t1) );
fim FAN_N3305_0 ( .fault(fault), .net(N3305), .FEN(FEN[1887]), .op(N3305_t0) );
fim FAN_N3305_1 ( .fault(fault), .net(N3305), .FEN(FEN[1888]), .op(N3305_t1) );
fim FAN_N3305_2 ( .fault(fault), .net(N3305), .FEN(FEN[1889]), .op(N3305_t2) );
fim FAN_N3314_0 ( .fault(fault), .net(N3314), .FEN(FEN[1890]), .op(N3314_t0) );
fim FAN_N3314_1 ( .fault(fault), .net(N3314), .FEN(FEN[1891]), .op(N3314_t1) );
fim FAN_N3311_0 ( .fault(fault), .net(N3311), .FEN(FEN[1892]), .op(N3311_t0) );
fim FAN_N3311_1 ( .fault(fault), .net(N3311), .FEN(FEN[1893]), .op(N3311_t1) );
fim FAN_N3317_0 ( .fault(fault), .net(N3317), .FEN(FEN[1894]), .op(N3317_t0) );
fim FAN_N3317_1 ( .fault(fault), .net(N3317), .FEN(FEN[1895]), .op(N3317_t1) );
fim FAN_N3317_2 ( .fault(fault), .net(N3317), .FEN(FEN[1896]), .op(N3317_t2) );
fim FAN_N3341_0 ( .fault(fault), .net(N3341), .FEN(FEN[1897]), .op(N3341_t0) );
fim FAN_N3341_1 ( .fault(fault), .net(N3341), .FEN(FEN[1898]), .op(N3341_t1) );
fim FAN_N996_0 ( .fault(fault), .net(N996), .FEN(FEN[1899]), .op(N996_t0) );
fim FAN_N996_1 ( .fault(fault), .net(N996), .FEN(FEN[1900]), .op(N996_t1) );
fim FAN_N3344_0 ( .fault(fault), .net(N3344), .FEN(FEN[1901]), .op(N3344_t0) );
fim FAN_N3344_1 ( .fault(fault), .net(N3344), .FEN(FEN[1902]), .op(N3344_t1) );
fim FAN_N3344_2 ( .fault(fault), .net(N3344), .FEN(FEN[1903]), .op(N3344_t2) );
fim FAN_N3353_0 ( .fault(fault), .net(N3353), .FEN(FEN[1904]), .op(N3353_t0) );
fim FAN_N3353_1 ( .fault(fault), .net(N3353), .FEN(FEN[1905]), .op(N3353_t1) );
fim FAN_N3350_0 ( .fault(fault), .net(N3350), .FEN(FEN[1906]), .op(N3350_t0) );
fim FAN_N3350_1 ( .fault(fault), .net(N3350), .FEN(FEN[1907]), .op(N3350_t1) );
fim FAN_N3356_0 ( .fault(fault), .net(N3356), .FEN(FEN[1908]), .op(N3356_t0) );
fim FAN_N3356_1 ( .fault(fault), .net(N3356), .FEN(FEN[1909]), .op(N3356_t1) );
fim FAN_N3356_2 ( .fault(fault), .net(N3356), .FEN(FEN[1910]), .op(N3356_t2) );
fim FAN_N3362_0 ( .fault(fault), .net(N3362), .FEN(FEN[1911]), .op(N3362_t0) );
fim FAN_N3362_1 ( .fault(fault), .net(N3362), .FEN(FEN[1912]), .op(N3362_t1) );
fim FAN_N1239_0 ( .fault(fault), .net(N1239), .FEN(FEN[1913]), .op(N1239_t0) );
fim FAN_N1239_1 ( .fault(fault), .net(N1239), .FEN(FEN[1914]), .op(N1239_t1) );
fim FAN_N3365_0 ( .fault(fault), .net(N3365), .FEN(FEN[1915]), .op(N3365_t0) );
fim FAN_N3365_1 ( .fault(fault), .net(N3365), .FEN(FEN[1916]), .op(N3365_t1) );
fim FAN_N564_0 ( .fault(fault), .net(N564), .FEN(FEN[1917]), .op(N564_t0) );
fim FAN_N564_1 ( .fault(fault), .net(N564), .FEN(FEN[1918]), .op(N564_t1) );
fim FAN_N3368_0 ( .fault(fault), .net(N3368), .FEN(FEN[1919]), .op(N3368_t0) );
fim FAN_N3368_1 ( .fault(fault), .net(N3368), .FEN(FEN[1920]), .op(N3368_t1) );
fim FAN_N612_0 ( .fault(fault), .net(N612), .FEN(FEN[1921]), .op(N612_t0) );
fim FAN_N612_1 ( .fault(fault), .net(N612), .FEN(FEN[1922]), .op(N612_t1) );
fim FAN_N3371_0 ( .fault(fault), .net(N3371), .FEN(FEN[1923]), .op(N3371_t0) );
fim FAN_N3371_1 ( .fault(fault), .net(N3371), .FEN(FEN[1924]), .op(N3371_t1) );
fim FAN_N660_0 ( .fault(fault), .net(N660), .FEN(FEN[1925]), .op(N660_t0) );
fim FAN_N660_1 ( .fault(fault), .net(N660), .FEN(FEN[1926]), .op(N660_t1) );
fim FAN_N3374_0 ( .fault(fault), .net(N3374), .FEN(FEN[1927]), .op(N3374_t0) );
fim FAN_N3374_1 ( .fault(fault), .net(N3374), .FEN(FEN[1928]), .op(N3374_t1) );
fim FAN_N708_0 ( .fault(fault), .net(N708), .FEN(FEN[1929]), .op(N708_t0) );
fim FAN_N708_1 ( .fault(fault), .net(N708), .FEN(FEN[1930]), .op(N708_t1) );
fim FAN_N3377_0 ( .fault(fault), .net(N3377), .FEN(FEN[1931]), .op(N3377_t0) );
fim FAN_N3377_1 ( .fault(fault), .net(N3377), .FEN(FEN[1932]), .op(N3377_t1) );
fim FAN_N756_0 ( .fault(fault), .net(N756), .FEN(FEN[1933]), .op(N756_t0) );
fim FAN_N756_1 ( .fault(fault), .net(N756), .FEN(FEN[1934]), .op(N756_t1) );
fim FAN_N3380_0 ( .fault(fault), .net(N3380), .FEN(FEN[1935]), .op(N3380_t0) );
fim FAN_N3380_1 ( .fault(fault), .net(N3380), .FEN(FEN[1936]), .op(N3380_t1) );
fim FAN_N804_0 ( .fault(fault), .net(N804), .FEN(FEN[1937]), .op(N804_t0) );
fim FAN_N804_1 ( .fault(fault), .net(N804), .FEN(FEN[1938]), .op(N804_t1) );
fim FAN_N3383_0 ( .fault(fault), .net(N3383), .FEN(FEN[1939]), .op(N3383_t0) );
fim FAN_N3383_1 ( .fault(fault), .net(N3383), .FEN(FEN[1940]), .op(N3383_t1) );
fim FAN_N852_0 ( .fault(fault), .net(N852), .FEN(FEN[1941]), .op(N852_t0) );
fim FAN_N852_1 ( .fault(fault), .net(N852), .FEN(FEN[1942]), .op(N852_t1) );
fim FAN_N3386_0 ( .fault(fault), .net(N3386), .FEN(FEN[1943]), .op(N3386_t0) );
fim FAN_N3386_1 ( .fault(fault), .net(N3386), .FEN(FEN[1944]), .op(N3386_t1) );
fim FAN_N900_0 ( .fault(fault), .net(N900), .FEN(FEN[1945]), .op(N900_t0) );
fim FAN_N900_1 ( .fault(fault), .net(N900), .FEN(FEN[1946]), .op(N900_t1) );
fim FAN_N3389_0 ( .fault(fault), .net(N3389), .FEN(FEN[1947]), .op(N3389_t0) );
fim FAN_N3389_1 ( .fault(fault), .net(N3389), .FEN(FEN[1948]), .op(N3389_t1) );
fim FAN_N948_0 ( .fault(fault), .net(N948), .FEN(FEN[1949]), .op(N948_t0) );
fim FAN_N948_1 ( .fault(fault), .net(N948), .FEN(FEN[1950]), .op(N948_t1) );
fim FAN_N3392_0 ( .fault(fault), .net(N3392), .FEN(FEN[1951]), .op(N3392_t0) );
fim FAN_N3392_1 ( .fault(fault), .net(N3392), .FEN(FEN[1952]), .op(N3392_t1) );
fim FAN_N3392_2 ( .fault(fault), .net(N3392), .FEN(FEN[1953]), .op(N3392_t2) );
fim FAN_N3401_0 ( .fault(fault), .net(N3401), .FEN(FEN[1954]), .op(N3401_t0) );
fim FAN_N3401_1 ( .fault(fault), .net(N3401), .FEN(FEN[1955]), .op(N3401_t1) );
fim FAN_N3398_0 ( .fault(fault), .net(N3398), .FEN(FEN[1956]), .op(N3398_t0) );
fim FAN_N3398_1 ( .fault(fault), .net(N3398), .FEN(FEN[1957]), .op(N3398_t1) );
fim FAN_N3404_0 ( .fault(fault), .net(N3404), .FEN(FEN[1958]), .op(N3404_t0) );
fim FAN_N3404_1 ( .fault(fault), .net(N3404), .FEN(FEN[1959]), .op(N3404_t1) );
fim FAN_N3404_2 ( .fault(fault), .net(N3404), .FEN(FEN[1960]), .op(N3404_t2) );
fim FAN_N3410_0 ( .fault(fault), .net(N3410), .FEN(FEN[1961]), .op(N3410_t0) );
fim FAN_N3410_1 ( .fault(fault), .net(N3410), .FEN(FEN[1962]), .op(N3410_t1) );
fim FAN_N1191_0 ( .fault(fault), .net(N1191), .FEN(FEN[1963]), .op(N1191_t0) );
fim FAN_N1191_1 ( .fault(fault), .net(N1191), .FEN(FEN[1964]), .op(N1191_t1) );
fim FAN_N3413_0 ( .fault(fault), .net(N3413), .FEN(FEN[1965]), .op(N3413_t0) );
fim FAN_N3413_1 ( .fault(fault), .net(N3413), .FEN(FEN[1966]), .op(N3413_t1) );
fim FAN_N3413_2 ( .fault(fault), .net(N3413), .FEN(FEN[1967]), .op(N3413_t2) );
fim FAN_N3417_0 ( .fault(fault), .net(N3417), .FEN(FEN[1968]), .op(N3417_t0) );
fim FAN_N3417_1 ( .fault(fault), .net(N3417), .FEN(FEN[1969]), .op(N3417_t1) );
fim FAN_N3417_2 ( .fault(fault), .net(N3417), .FEN(FEN[1970]), .op(N3417_t2) );
fim FAN_N3421_0 ( .fault(fault), .net(N3421), .FEN(FEN[1971]), .op(N3421_t0) );
fim FAN_N3421_1 ( .fault(fault), .net(N3421), .FEN(FEN[1972]), .op(N3421_t1) );
fim FAN_N3421_2 ( .fault(fault), .net(N3421), .FEN(FEN[1973]), .op(N3421_t2) );
fim FAN_N3425_0 ( .fault(fault), .net(N3425), .FEN(FEN[1974]), .op(N3425_t0) );
fim FAN_N3425_1 ( .fault(fault), .net(N3425), .FEN(FEN[1975]), .op(N3425_t1) );
fim FAN_N3425_2 ( .fault(fault), .net(N3425), .FEN(FEN[1976]), .op(N3425_t2) );
fim FAN_N3429_0 ( .fault(fault), .net(N3429), .FEN(FEN[1977]), .op(N3429_t0) );
fim FAN_N3429_1 ( .fault(fault), .net(N3429), .FEN(FEN[1978]), .op(N3429_t1) );
fim FAN_N3429_2 ( .fault(fault), .net(N3429), .FEN(FEN[1979]), .op(N3429_t2) );
fim FAN_N3433_0 ( .fault(fault), .net(N3433), .FEN(FEN[1980]), .op(N3433_t0) );
fim FAN_N3433_1 ( .fault(fault), .net(N3433), .FEN(FEN[1981]), .op(N3433_t1) );
fim FAN_N3433_2 ( .fault(fault), .net(N3433), .FEN(FEN[1982]), .op(N3433_t2) );
fim FAN_N3437_0 ( .fault(fault), .net(N3437), .FEN(FEN[1983]), .op(N3437_t0) );
fim FAN_N3437_1 ( .fault(fault), .net(N3437), .FEN(FEN[1984]), .op(N3437_t1) );
fim FAN_N3437_2 ( .fault(fault), .net(N3437), .FEN(FEN[1985]), .op(N3437_t2) );
fim FAN_N3441_0 ( .fault(fault), .net(N3441), .FEN(FEN[1986]), .op(N3441_t0) );
fim FAN_N3441_1 ( .fault(fault), .net(N3441), .FEN(FEN[1987]), .op(N3441_t1) );
fim FAN_N3441_2 ( .fault(fault), .net(N3441), .FEN(FEN[1988]), .op(N3441_t2) );
fim FAN_N3445_0 ( .fault(fault), .net(N3445), .FEN(FEN[1989]), .op(N3445_t0) );
fim FAN_N3445_1 ( .fault(fault), .net(N3445), .FEN(FEN[1990]), .op(N3445_t1) );
fim FAN_N3445_2 ( .fault(fault), .net(N3445), .FEN(FEN[1991]), .op(N3445_t2) );
fim FAN_N3449_0 ( .fault(fault), .net(N3449), .FEN(FEN[1992]), .op(N3449_t0) );
fim FAN_N3449_1 ( .fault(fault), .net(N3449), .FEN(FEN[1993]), .op(N3449_t1) );
fim FAN_N3449_2 ( .fault(fault), .net(N3449), .FEN(FEN[1994]), .op(N3449_t2) );
fim FAN_N3458_0 ( .fault(fault), .net(N3458), .FEN(FEN[1995]), .op(N3458_t0) );
fim FAN_N3458_1 ( .fault(fault), .net(N3458), .FEN(FEN[1996]), .op(N3458_t1) );
fim FAN_N3455_0 ( .fault(fault), .net(N3455), .FEN(FEN[1997]), .op(N3455_t0) );
fim FAN_N3455_1 ( .fault(fault), .net(N3455), .FEN(FEN[1998]), .op(N3455_t1) );
fim FAN_N3461_0 ( .fault(fault), .net(N3461), .FEN(FEN[1999]), .op(N3461_t0) );
fim FAN_N3461_1 ( .fault(fault), .net(N3461), .FEN(FEN[2000]), .op(N3461_t1) );
fim FAN_N3461_2 ( .fault(fault), .net(N3461), .FEN(FEN[2001]), .op(N3461_t2) );
fim FAN_N3467_0 ( .fault(fault), .net(N3467), .FEN(FEN[2002]), .op(N3467_t0) );
fim FAN_N3467_1 ( .fault(fault), .net(N3467), .FEN(FEN[2003]), .op(N3467_t1) );
fim FAN_N1143_0 ( .fault(fault), .net(N1143), .FEN(FEN[2004]), .op(N1143_t0) );
fim FAN_N1143_1 ( .fault(fault), .net(N1143), .FEN(FEN[2005]), .op(N1143_t1) );
fim FAN_N3470_0 ( .fault(fault), .net(N3470), .FEN(FEN[2006]), .op(N3470_t0) );
fim FAN_N3470_1 ( .fault(fault), .net(N3470), .FEN(FEN[2007]), .op(N3470_t1) );
fim FAN_N3470_2 ( .fault(fault), .net(N3470), .FEN(FEN[2008]), .op(N3470_t2) );
fim FAN_N1287_0 ( .fault(fault), .net(N1287), .FEN(FEN[2009]), .op(N1287_t0) );
fim FAN_N1287_1 ( .fault(fault), .net(N1287), .FEN(FEN[2010]), .op(N1287_t1) );
fim FAN_N3476_0 ( .fault(fault), .net(N3476), .FEN(FEN[2011]), .op(N3476_t0) );
fim FAN_N3476_1 ( .fault(fault), .net(N3476), .FEN(FEN[2012]), .op(N3476_t1) );
fim FAN_N3524_0 ( .fault(fault), .net(N3524), .FEN(FEN[2013]), .op(N3524_t0) );
fim FAN_N3524_1 ( .fault(fault), .net(N3524), .FEN(FEN[2014]), .op(N3524_t1) );
fim FAN_N3521_0 ( .fault(fault), .net(N3521), .FEN(FEN[2015]), .op(N3521_t0) );
fim FAN_N3521_1 ( .fault(fault), .net(N3521), .FEN(FEN[2016]), .op(N3521_t1) );
fim FAN_N3527_0 ( .fault(fault), .net(N3527), .FEN(FEN[2017]), .op(N3527_t0) );
fim FAN_N3527_1 ( .fault(fault), .net(N3527), .FEN(FEN[2018]), .op(N3527_t1) );
fim FAN_N3527_2 ( .fault(fault), .net(N3527), .FEN(FEN[2019]), .op(N3527_t2) );
fim FAN_N3533_0 ( .fault(fault), .net(N3533), .FEN(FEN[2020]), .op(N3533_t0) );
fim FAN_N3533_1 ( .fault(fault), .net(N3533), .FEN(FEN[2021]), .op(N3533_t1) );
fim FAN_N1095_0 ( .fault(fault), .net(N1095), .FEN(FEN[2022]), .op(N1095_t0) );
fim FAN_N1095_1 ( .fault(fault), .net(N1095), .FEN(FEN[2023]), .op(N1095_t1) );
fim FAN_N3536_0 ( .fault(fault), .net(N3536), .FEN(FEN[2024]), .op(N3536_t0) );
fim FAN_N3536_1 ( .fault(fault), .net(N3536), .FEN(FEN[2025]), .op(N3536_t1) );
fim FAN_N3536_2 ( .fault(fault), .net(N3536), .FEN(FEN[2026]), .op(N3536_t2) );
fim FAN_N3545_0 ( .fault(fault), .net(N3545), .FEN(FEN[2027]), .op(N3545_t0) );
fim FAN_N3545_1 ( .fault(fault), .net(N3545), .FEN(FEN[2028]), .op(N3545_t1) );
fim FAN_N3542_0 ( .fault(fault), .net(N3542), .FEN(FEN[2029]), .op(N3542_t0) );
fim FAN_N3542_1 ( .fault(fault), .net(N3542), .FEN(FEN[2030]), .op(N3542_t1) );
fim FAN_N3548_0 ( .fault(fault), .net(N3548), .FEN(FEN[2031]), .op(N3548_t0) );
fim FAN_N3548_1 ( .fault(fault), .net(N3548), .FEN(FEN[2032]), .op(N3548_t1) );
fim FAN_N3548_2 ( .fault(fault), .net(N3548), .FEN(FEN[2033]), .op(N3548_t2) );
fim FAN_N3553_0 ( .fault(fault), .net(N3553), .FEN(FEN[2034]), .op(N3553_t0) );
fim FAN_N3553_1 ( .fault(fault), .net(N3553), .FEN(FEN[2035]), .op(N3553_t1) );
fim FAN_N3481_0 ( .fault(fault), .net(N3481), .FEN(FEN[2036]), .op(N3481_t0) );
fim FAN_N3481_1 ( .fault(fault), .net(N3481), .FEN(FEN[2037]), .op(N3481_t1) );
fim FAN_N3556_0 ( .fault(fault), .net(N3556), .FEN(FEN[2038]), .op(N3556_t0) );
fim FAN_N3556_1 ( .fault(fault), .net(N3556), .FEN(FEN[2039]), .op(N3556_t1) );
fim FAN_N3486_0 ( .fault(fault), .net(N3486), .FEN(FEN[2040]), .op(N3486_t0) );
fim FAN_N3486_1 ( .fault(fault), .net(N3486), .FEN(FEN[2041]), .op(N3486_t1) );
fim FAN_N3559_0 ( .fault(fault), .net(N3559), .FEN(FEN[2042]), .op(N3559_t0) );
fim FAN_N3559_1 ( .fault(fault), .net(N3559), .FEN(FEN[2043]), .op(N3559_t1) );
fim FAN_N3491_0 ( .fault(fault), .net(N3491), .FEN(FEN[2044]), .op(N3491_t0) );
fim FAN_N3491_1 ( .fault(fault), .net(N3491), .FEN(FEN[2045]), .op(N3491_t1) );
fim FAN_N3562_0 ( .fault(fault), .net(N3562), .FEN(FEN[2046]), .op(N3562_t0) );
fim FAN_N3562_1 ( .fault(fault), .net(N3562), .FEN(FEN[2047]), .op(N3562_t1) );
fim FAN_N3496_0 ( .fault(fault), .net(N3496), .FEN(FEN[2048]), .op(N3496_t0) );
fim FAN_N3496_1 ( .fault(fault), .net(N3496), .FEN(FEN[2049]), .op(N3496_t1) );
fim FAN_N3565_0 ( .fault(fault), .net(N3565), .FEN(FEN[2050]), .op(N3565_t0) );
fim FAN_N3565_1 ( .fault(fault), .net(N3565), .FEN(FEN[2051]), .op(N3565_t1) );
fim FAN_N3501_0 ( .fault(fault), .net(N3501), .FEN(FEN[2052]), .op(N3501_t0) );
fim FAN_N3501_1 ( .fault(fault), .net(N3501), .FEN(FEN[2053]), .op(N3501_t1) );
fim FAN_N3568_0 ( .fault(fault), .net(N3568), .FEN(FEN[2054]), .op(N3568_t0) );
fim FAN_N3568_1 ( .fault(fault), .net(N3568), .FEN(FEN[2055]), .op(N3568_t1) );
fim FAN_N3506_0 ( .fault(fault), .net(N3506), .FEN(FEN[2056]), .op(N3506_t0) );
fim FAN_N3506_1 ( .fault(fault), .net(N3506), .FEN(FEN[2057]), .op(N3506_t1) );
fim FAN_N3571_0 ( .fault(fault), .net(N3571), .FEN(FEN[2058]), .op(N3571_t0) );
fim FAN_N3571_1 ( .fault(fault), .net(N3571), .FEN(FEN[2059]), .op(N3571_t1) );
fim FAN_N3511_0 ( .fault(fault), .net(N3511), .FEN(FEN[2060]), .op(N3511_t0) );
fim FAN_N3511_1 ( .fault(fault), .net(N3511), .FEN(FEN[2061]), .op(N3511_t1) );
fim FAN_N3574_0 ( .fault(fault), .net(N3574), .FEN(FEN[2062]), .op(N3574_t0) );
fim FAN_N3574_1 ( .fault(fault), .net(N3574), .FEN(FEN[2063]), .op(N3574_t1) );
fim FAN_N3516_0 ( .fault(fault), .net(N3516), .FEN(FEN[2064]), .op(N3516_t0) );
fim FAN_N3516_1 ( .fault(fault), .net(N3516), .FEN(FEN[2065]), .op(N3516_t1) );
fim FAN_N3577_0 ( .fault(fault), .net(N3577), .FEN(FEN[2066]), .op(N3577_t0) );
fim FAN_N3577_1 ( .fault(fault), .net(N3577), .FEN(FEN[2067]), .op(N3577_t1) );
fim FAN_N3577_2 ( .fault(fault), .net(N3577), .FEN(FEN[2068]), .op(N3577_t2) );
fim FAN_N3583_0 ( .fault(fault), .net(N3583), .FEN(FEN[2069]), .op(N3583_t0) );
fim FAN_N3583_1 ( .fault(fault), .net(N3583), .FEN(FEN[2070]), .op(N3583_t1) );
fim FAN_N1047_0 ( .fault(fault), .net(N1047), .FEN(FEN[2071]), .op(N1047_t0) );
fim FAN_N1047_1 ( .fault(fault), .net(N1047), .FEN(FEN[2072]), .op(N1047_t1) );
fim FAN_N3586_0 ( .fault(fault), .net(N3586), .FEN(FEN[2073]), .op(N3586_t0) );
fim FAN_N3586_1 ( .fault(fault), .net(N3586), .FEN(FEN[2074]), .op(N3586_t1) );
fim FAN_N3586_2 ( .fault(fault), .net(N3586), .FEN(FEN[2075]), .op(N3586_t2) );
fim FAN_N3595_0 ( .fault(fault), .net(N3595), .FEN(FEN[2076]), .op(N3595_t0) );
fim FAN_N3595_1 ( .fault(fault), .net(N3595), .FEN(FEN[2077]), .op(N3595_t1) );
fim FAN_N3592_0 ( .fault(fault), .net(N3592), .FEN(FEN[2078]), .op(N3592_t0) );
fim FAN_N3592_1 ( .fault(fault), .net(N3592), .FEN(FEN[2079]), .op(N3592_t1) );
fim FAN_N3598_0 ( .fault(fault), .net(N3598), .FEN(FEN[2080]), .op(N3598_t0) );
fim FAN_N3598_1 ( .fault(fault), .net(N3598), .FEN(FEN[2081]), .op(N3598_t1) );
fim FAN_N3598_2 ( .fault(fault), .net(N3598), .FEN(FEN[2082]), .op(N3598_t2) );
fim FAN_N3604_0 ( .fault(fault), .net(N3604), .FEN(FEN[2083]), .op(N3604_t0) );
fim FAN_N3604_1 ( .fault(fault), .net(N3604), .FEN(FEN[2084]), .op(N3604_t1) );
fim FAN_N3604_2 ( .fault(fault), .net(N3604), .FEN(FEN[2085]), .op(N3604_t2) );
fim FAN_N3608_0 ( .fault(fault), .net(N3608), .FEN(FEN[2086]), .op(N3608_t0) );
fim FAN_N3608_1 ( .fault(fault), .net(N3608), .FEN(FEN[2087]), .op(N3608_t1) );
fim FAN_N3608_2 ( .fault(fault), .net(N3608), .FEN(FEN[2088]), .op(N3608_t2) );
fim FAN_N3612_0 ( .fault(fault), .net(N3612), .FEN(FEN[2089]), .op(N3612_t0) );
fim FAN_N3612_1 ( .fault(fault), .net(N3612), .FEN(FEN[2090]), .op(N3612_t1) );
fim FAN_N3612_2 ( .fault(fault), .net(N3612), .FEN(FEN[2091]), .op(N3612_t2) );
fim FAN_N3616_0 ( .fault(fault), .net(N3616), .FEN(FEN[2092]), .op(N3616_t0) );
fim FAN_N3616_1 ( .fault(fault), .net(N3616), .FEN(FEN[2093]), .op(N3616_t1) );
fim FAN_N3616_2 ( .fault(fault), .net(N3616), .FEN(FEN[2094]), .op(N3616_t2) );
fim FAN_N3620_0 ( .fault(fault), .net(N3620), .FEN(FEN[2095]), .op(N3620_t0) );
fim FAN_N3620_1 ( .fault(fault), .net(N3620), .FEN(FEN[2096]), .op(N3620_t1) );
fim FAN_N3620_2 ( .fault(fault), .net(N3620), .FEN(FEN[2097]), .op(N3620_t2) );
fim FAN_N3624_0 ( .fault(fault), .net(N3624), .FEN(FEN[2098]), .op(N3624_t0) );
fim FAN_N3624_1 ( .fault(fault), .net(N3624), .FEN(FEN[2099]), .op(N3624_t1) );
fim FAN_N3624_2 ( .fault(fault), .net(N3624), .FEN(FEN[2100]), .op(N3624_t2) );
fim FAN_N3628_0 ( .fault(fault), .net(N3628), .FEN(FEN[2101]), .op(N3628_t0) );
fim FAN_N3628_1 ( .fault(fault), .net(N3628), .FEN(FEN[2102]), .op(N3628_t1) );
fim FAN_N3628_2 ( .fault(fault), .net(N3628), .FEN(FEN[2103]), .op(N3628_t2) );
fim FAN_N3632_0 ( .fault(fault), .net(N3632), .FEN(FEN[2104]), .op(N3632_t0) );
fim FAN_N3632_1 ( .fault(fault), .net(N3632), .FEN(FEN[2105]), .op(N3632_t1) );
fim FAN_N3632_2 ( .fault(fault), .net(N3632), .FEN(FEN[2106]), .op(N3632_t2) );
fim FAN_N3638_0 ( .fault(fault), .net(N3638), .FEN(FEN[2107]), .op(N3638_t0) );
fim FAN_N3638_1 ( .fault(fault), .net(N3638), .FEN(FEN[2108]), .op(N3638_t1) );
fim FAN_N999_0 ( .fault(fault), .net(N999), .FEN(FEN[2109]), .op(N999_t0) );
fim FAN_N999_1 ( .fault(fault), .net(N999), .FEN(FEN[2110]), .op(N999_t1) );
fim FAN_N3641_0 ( .fault(fault), .net(N3641), .FEN(FEN[2111]), .op(N3641_t0) );
fim FAN_N3641_1 ( .fault(fault), .net(N3641), .FEN(FEN[2112]), .op(N3641_t1) );
fim FAN_N3641_2 ( .fault(fault), .net(N3641), .FEN(FEN[2113]), .op(N3641_t2) );
fim FAN_N3650_0 ( .fault(fault), .net(N3650), .FEN(FEN[2114]), .op(N3650_t0) );
fim FAN_N3650_1 ( .fault(fault), .net(N3650), .FEN(FEN[2115]), .op(N3650_t1) );
fim FAN_N3647_0 ( .fault(fault), .net(N3647), .FEN(FEN[2116]), .op(N3647_t0) );
fim FAN_N3647_1 ( .fault(fault), .net(N3647), .FEN(FEN[2117]), .op(N3647_t1) );
fim FAN_N3653_0 ( .fault(fault), .net(N3653), .FEN(FEN[2118]), .op(N3653_t0) );
fim FAN_N3653_1 ( .fault(fault), .net(N3653), .FEN(FEN[2119]), .op(N3653_t1) );
fim FAN_N3653_2 ( .fault(fault), .net(N3653), .FEN(FEN[2120]), .op(N3653_t2) );
fim FAN_N3659_0 ( .fault(fault), .net(N3659), .FEN(FEN[2121]), .op(N3659_t0) );
fim FAN_N3659_1 ( .fault(fault), .net(N3659), .FEN(FEN[2122]), .op(N3659_t1) );
fim FAN_N1242_0 ( .fault(fault), .net(N1242), .FEN(FEN[2123]), .op(N1242_t0) );
fim FAN_N1242_1 ( .fault(fault), .net(N1242), .FEN(FEN[2124]), .op(N1242_t1) );
fim FAN_N3678_0 ( .fault(fault), .net(N3678), .FEN(FEN[2125]), .op(N3678_t0) );
fim FAN_N3678_1 ( .fault(fault), .net(N3678), .FEN(FEN[2126]), .op(N3678_t1) );
fim FAN_N951_0 ( .fault(fault), .net(N951), .FEN(FEN[2127]), .op(N951_t0) );
fim FAN_N951_1 ( .fault(fault), .net(N951), .FEN(FEN[2128]), .op(N951_t1) );
fim FAN_N3681_0 ( .fault(fault), .net(N3681), .FEN(FEN[2129]), .op(N3681_t0) );
fim FAN_N3681_1 ( .fault(fault), .net(N3681), .FEN(FEN[2130]), .op(N3681_t1) );
fim FAN_N3681_2 ( .fault(fault), .net(N3681), .FEN(FEN[2131]), .op(N3681_t2) );
fim FAN_N3690_0 ( .fault(fault), .net(N3690), .FEN(FEN[2132]), .op(N3690_t0) );
fim FAN_N3690_1 ( .fault(fault), .net(N3690), .FEN(FEN[2133]), .op(N3690_t1) );
fim FAN_N3687_0 ( .fault(fault), .net(N3687), .FEN(FEN[2134]), .op(N3687_t0) );
fim FAN_N3687_1 ( .fault(fault), .net(N3687), .FEN(FEN[2135]), .op(N3687_t1) );
fim FAN_N3693_0 ( .fault(fault), .net(N3693), .FEN(FEN[2136]), .op(N3693_t0) );
fim FAN_N3693_1 ( .fault(fault), .net(N3693), .FEN(FEN[2137]), .op(N3693_t1) );
fim FAN_N3693_2 ( .fault(fault), .net(N3693), .FEN(FEN[2138]), .op(N3693_t2) );
fim FAN_N3699_0 ( .fault(fault), .net(N3699), .FEN(FEN[2139]), .op(N3699_t0) );
fim FAN_N3699_1 ( .fault(fault), .net(N3699), .FEN(FEN[2140]), .op(N3699_t1) );
fim FAN_N1194_0 ( .fault(fault), .net(N1194), .FEN(FEN[2141]), .op(N1194_t0) );
fim FAN_N1194_1 ( .fault(fault), .net(N1194), .FEN(FEN[2142]), .op(N1194_t1) );
fim FAN_N3702_0 ( .fault(fault), .net(N3702), .FEN(FEN[2143]), .op(N3702_t0) );
fim FAN_N3702_1 ( .fault(fault), .net(N3702), .FEN(FEN[2144]), .op(N3702_t1) );
fim FAN_N3702_2 ( .fault(fault), .net(N3702), .FEN(FEN[2145]), .op(N3702_t2) );
fim FAN_N3706_0 ( .fault(fault), .net(N3706), .FEN(FEN[2146]), .op(N3706_t0) );
fim FAN_N3706_1 ( .fault(fault), .net(N3706), .FEN(FEN[2147]), .op(N3706_t1) );
fim FAN_N567_0 ( .fault(fault), .net(N567), .FEN(FEN[2148]), .op(N567_t0) );
fim FAN_N567_1 ( .fault(fault), .net(N567), .FEN(FEN[2149]), .op(N567_t1) );
fim FAN_N3709_0 ( .fault(fault), .net(N3709), .FEN(FEN[2150]), .op(N3709_t0) );
fim FAN_N3709_1 ( .fault(fault), .net(N3709), .FEN(FEN[2151]), .op(N3709_t1) );
fim FAN_N615_0 ( .fault(fault), .net(N615), .FEN(FEN[2152]), .op(N615_t0) );
fim FAN_N615_1 ( .fault(fault), .net(N615), .FEN(FEN[2153]), .op(N615_t1) );
fim FAN_N3712_0 ( .fault(fault), .net(N3712), .FEN(FEN[2154]), .op(N3712_t0) );
fim FAN_N3712_1 ( .fault(fault), .net(N3712), .FEN(FEN[2155]), .op(N3712_t1) );
fim FAN_N663_0 ( .fault(fault), .net(N663), .FEN(FEN[2156]), .op(N663_t0) );
fim FAN_N663_1 ( .fault(fault), .net(N663), .FEN(FEN[2157]), .op(N663_t1) );
fim FAN_N3715_0 ( .fault(fault), .net(N3715), .FEN(FEN[2158]), .op(N3715_t0) );
fim FAN_N3715_1 ( .fault(fault), .net(N3715), .FEN(FEN[2159]), .op(N3715_t1) );
fim FAN_N711_0 ( .fault(fault), .net(N711), .FEN(FEN[2160]), .op(N711_t0) );
fim FAN_N711_1 ( .fault(fault), .net(N711), .FEN(FEN[2161]), .op(N711_t1) );
fim FAN_N3718_0 ( .fault(fault), .net(N3718), .FEN(FEN[2162]), .op(N3718_t0) );
fim FAN_N3718_1 ( .fault(fault), .net(N3718), .FEN(FEN[2163]), .op(N3718_t1) );
fim FAN_N759_0 ( .fault(fault), .net(N759), .FEN(FEN[2164]), .op(N759_t0) );
fim FAN_N759_1 ( .fault(fault), .net(N759), .FEN(FEN[2165]), .op(N759_t1) );
fim FAN_N3721_0 ( .fault(fault), .net(N3721), .FEN(FEN[2166]), .op(N3721_t0) );
fim FAN_N3721_1 ( .fault(fault), .net(N3721), .FEN(FEN[2167]), .op(N3721_t1) );
fim FAN_N807_0 ( .fault(fault), .net(N807), .FEN(FEN[2168]), .op(N807_t0) );
fim FAN_N807_1 ( .fault(fault), .net(N807), .FEN(FEN[2169]), .op(N807_t1) );
fim FAN_N3724_0 ( .fault(fault), .net(N3724), .FEN(FEN[2170]), .op(N3724_t0) );
fim FAN_N3724_1 ( .fault(fault), .net(N3724), .FEN(FEN[2171]), .op(N3724_t1) );
fim FAN_N855_0 ( .fault(fault), .net(N855), .FEN(FEN[2172]), .op(N855_t0) );
fim FAN_N855_1 ( .fault(fault), .net(N855), .FEN(FEN[2173]), .op(N855_t1) );
fim FAN_N3727_0 ( .fault(fault), .net(N3727), .FEN(FEN[2174]), .op(N3727_t0) );
fim FAN_N3727_1 ( .fault(fault), .net(N3727), .FEN(FEN[2175]), .op(N3727_t1) );
fim FAN_N903_0 ( .fault(fault), .net(N903), .FEN(FEN[2176]), .op(N903_t0) );
fim FAN_N903_1 ( .fault(fault), .net(N903), .FEN(FEN[2177]), .op(N903_t1) );
fim FAN_N3730_0 ( .fault(fault), .net(N3730), .FEN(FEN[2178]), .op(N3730_t0) );
fim FAN_N3730_1 ( .fault(fault), .net(N3730), .FEN(FEN[2179]), .op(N3730_t1) );
fim FAN_N3730_2 ( .fault(fault), .net(N3730), .FEN(FEN[2180]), .op(N3730_t2) );
fim FAN_N3739_0 ( .fault(fault), .net(N3739), .FEN(FEN[2181]), .op(N3739_t0) );
fim FAN_N3739_1 ( .fault(fault), .net(N3739), .FEN(FEN[2182]), .op(N3739_t1) );
fim FAN_N3736_0 ( .fault(fault), .net(N3736), .FEN(FEN[2183]), .op(N3736_t0) );
fim FAN_N3736_1 ( .fault(fault), .net(N3736), .FEN(FEN[2184]), .op(N3736_t1) );
fim FAN_N3742_0 ( .fault(fault), .net(N3742), .FEN(FEN[2185]), .op(N3742_t0) );
fim FAN_N3742_1 ( .fault(fault), .net(N3742), .FEN(FEN[2186]), .op(N3742_t1) );
fim FAN_N3742_2 ( .fault(fault), .net(N3742), .FEN(FEN[2187]), .op(N3742_t2) );
fim FAN_N3748_0 ( .fault(fault), .net(N3748), .FEN(FEN[2188]), .op(N3748_t0) );
fim FAN_N3748_1 ( .fault(fault), .net(N3748), .FEN(FEN[2189]), .op(N3748_t1) );
fim FAN_N1146_0 ( .fault(fault), .net(N1146), .FEN(FEN[2190]), .op(N1146_t0) );
fim FAN_N1146_1 ( .fault(fault), .net(N1146), .FEN(FEN[2191]), .op(N1146_t1) );
fim FAN_N3751_0 ( .fault(fault), .net(N3751), .FEN(FEN[2192]), .op(N3751_t0) );
fim FAN_N3751_1 ( .fault(fault), .net(N3751), .FEN(FEN[2193]), .op(N3751_t1) );
fim FAN_N3751_2 ( .fault(fault), .net(N3751), .FEN(FEN[2194]), .op(N3751_t2) );
fim FAN_N1290_0 ( .fault(fault), .net(N1290), .FEN(FEN[2195]), .op(N1290_t0) );
fim FAN_N1290_1 ( .fault(fault), .net(N1290), .FEN(FEN[2196]), .op(N1290_t1) );
fim FAN_N3757_0 ( .fault(fault), .net(N3757), .FEN(FEN[2197]), .op(N3757_t0) );
fim FAN_N3757_1 ( .fault(fault), .net(N3757), .FEN(FEN[2198]), .op(N3757_t1) );
fim FAN_N3760_0 ( .fault(fault), .net(N3760), .FEN(FEN[2199]), .op(N3760_t0) );
fim FAN_N3760_1 ( .fault(fault), .net(N3760), .FEN(FEN[2200]), .op(N3760_t1) );
fim FAN_N3760_2 ( .fault(fault), .net(N3760), .FEN(FEN[2201]), .op(N3760_t2) );
fim FAN_N3764_0 ( .fault(fault), .net(N3764), .FEN(FEN[2202]), .op(N3764_t0) );
fim FAN_N3764_1 ( .fault(fault), .net(N3764), .FEN(FEN[2203]), .op(N3764_t1) );
fim FAN_N3764_2 ( .fault(fault), .net(N3764), .FEN(FEN[2204]), .op(N3764_t2) );
fim FAN_N3768_0 ( .fault(fault), .net(N3768), .FEN(FEN[2205]), .op(N3768_t0) );
fim FAN_N3768_1 ( .fault(fault), .net(N3768), .FEN(FEN[2206]), .op(N3768_t1) );
fim FAN_N3768_2 ( .fault(fault), .net(N3768), .FEN(FEN[2207]), .op(N3768_t2) );
fim FAN_N3772_0 ( .fault(fault), .net(N3772), .FEN(FEN[2208]), .op(N3772_t0) );
fim FAN_N3772_1 ( .fault(fault), .net(N3772), .FEN(FEN[2209]), .op(N3772_t1) );
fim FAN_N3772_2 ( .fault(fault), .net(N3772), .FEN(FEN[2210]), .op(N3772_t2) );
fim FAN_N3776_0 ( .fault(fault), .net(N3776), .FEN(FEN[2211]), .op(N3776_t0) );
fim FAN_N3776_1 ( .fault(fault), .net(N3776), .FEN(FEN[2212]), .op(N3776_t1) );
fim FAN_N3776_2 ( .fault(fault), .net(N3776), .FEN(FEN[2213]), .op(N3776_t2) );
fim FAN_N3780_0 ( .fault(fault), .net(N3780), .FEN(FEN[2214]), .op(N3780_t0) );
fim FAN_N3780_1 ( .fault(fault), .net(N3780), .FEN(FEN[2215]), .op(N3780_t1) );
fim FAN_N3780_2 ( .fault(fault), .net(N3780), .FEN(FEN[2216]), .op(N3780_t2) );
fim FAN_N3784_0 ( .fault(fault), .net(N3784), .FEN(FEN[2217]), .op(N3784_t0) );
fim FAN_N3784_1 ( .fault(fault), .net(N3784), .FEN(FEN[2218]), .op(N3784_t1) );
fim FAN_N3784_2 ( .fault(fault), .net(N3784), .FEN(FEN[2219]), .op(N3784_t2) );
fim FAN_N3788_0 ( .fault(fault), .net(N3788), .FEN(FEN[2220]), .op(N3788_t0) );
fim FAN_N3788_1 ( .fault(fault), .net(N3788), .FEN(FEN[2221]), .op(N3788_t1) );
fim FAN_N3788_2 ( .fault(fault), .net(N3788), .FEN(FEN[2222]), .op(N3788_t2) );
fim FAN_N3797_0 ( .fault(fault), .net(N3797), .FEN(FEN[2223]), .op(N3797_t0) );
fim FAN_N3797_1 ( .fault(fault), .net(N3797), .FEN(FEN[2224]), .op(N3797_t1) );
fim FAN_N3794_0 ( .fault(fault), .net(N3794), .FEN(FEN[2225]), .op(N3794_t0) );
fim FAN_N3794_1 ( .fault(fault), .net(N3794), .FEN(FEN[2226]), .op(N3794_t1) );
fim FAN_N3800_0 ( .fault(fault), .net(N3800), .FEN(FEN[2227]), .op(N3800_t0) );
fim FAN_N3800_1 ( .fault(fault), .net(N3800), .FEN(FEN[2228]), .op(N3800_t1) );
fim FAN_N3800_2 ( .fault(fault), .net(N3800), .FEN(FEN[2229]), .op(N3800_t2) );
fim FAN_N3806_0 ( .fault(fault), .net(N3806), .FEN(FEN[2230]), .op(N3806_t0) );
fim FAN_N3806_1 ( .fault(fault), .net(N3806), .FEN(FEN[2231]), .op(N3806_t1) );
fim FAN_N1098_0 ( .fault(fault), .net(N1098), .FEN(FEN[2232]), .op(N1098_t0) );
fim FAN_N1098_1 ( .fault(fault), .net(N1098), .FEN(FEN[2233]), .op(N1098_t1) );
fim FAN_N3809_0 ( .fault(fault), .net(N3809), .FEN(FEN[2234]), .op(N3809_t0) );
fim FAN_N3809_1 ( .fault(fault), .net(N3809), .FEN(FEN[2235]), .op(N3809_t1) );
fim FAN_N3809_2 ( .fault(fault), .net(N3809), .FEN(FEN[2236]), .op(N3809_t2) );
fim FAN_N3818_0 ( .fault(fault), .net(N3818), .FEN(FEN[2237]), .op(N3818_t0) );
fim FAN_N3818_1 ( .fault(fault), .net(N3818), .FEN(FEN[2238]), .op(N3818_t1) );
fim FAN_N3815_0 ( .fault(fault), .net(N3815), .FEN(FEN[2239]), .op(N3815_t0) );
fim FAN_N3815_1 ( .fault(fault), .net(N3815), .FEN(FEN[2240]), .op(N3815_t1) );
fim FAN_N3821_0 ( .fault(fault), .net(N3821), .FEN(FEN[2241]), .op(N3821_t0) );
fim FAN_N3821_1 ( .fault(fault), .net(N3821), .FEN(FEN[2242]), .op(N3821_t1) );
fim FAN_N3821_2 ( .fault(fault), .net(N3821), .FEN(FEN[2243]), .op(N3821_t2) );
fim FAN_N3865_0 ( .fault(fault), .net(N3865), .FEN(FEN[2244]), .op(N3865_t0) );
fim FAN_N3865_1 ( .fault(fault), .net(N3865), .FEN(FEN[2245]), .op(N3865_t1) );
fim FAN_N3862_0 ( .fault(fault), .net(N3862), .FEN(FEN[2246]), .op(N3862_t0) );
fim FAN_N3862_1 ( .fault(fault), .net(N3862), .FEN(FEN[2247]), .op(N3862_t1) );
fim FAN_N3868_0 ( .fault(fault), .net(N3868), .FEN(FEN[2248]), .op(N3868_t0) );
fim FAN_N3868_1 ( .fault(fault), .net(N3868), .FEN(FEN[2249]), .op(N3868_t1) );
fim FAN_N3868_2 ( .fault(fault), .net(N3868), .FEN(FEN[2250]), .op(N3868_t2) );
fim FAN_N3874_0 ( .fault(fault), .net(N3874), .FEN(FEN[2251]), .op(N3874_t0) );
fim FAN_N3874_1 ( .fault(fault), .net(N3874), .FEN(FEN[2252]), .op(N3874_t1) );
fim FAN_N1050_0 ( .fault(fault), .net(N1050), .FEN(FEN[2253]), .op(N1050_t0) );
fim FAN_N1050_1 ( .fault(fault), .net(N1050), .FEN(FEN[2254]), .op(N1050_t1) );
fim FAN_N3877_0 ( .fault(fault), .net(N3877), .FEN(FEN[2255]), .op(N3877_t0) );
fim FAN_N3877_1 ( .fault(fault), .net(N3877), .FEN(FEN[2256]), .op(N3877_t1) );
fim FAN_N3877_2 ( .fault(fault), .net(N3877), .FEN(FEN[2257]), .op(N3877_t2) );
fim FAN_N3886_0 ( .fault(fault), .net(N3886), .FEN(FEN[2258]), .op(N3886_t0) );
fim FAN_N3886_1 ( .fault(fault), .net(N3886), .FEN(FEN[2259]), .op(N3886_t1) );
fim FAN_N3883_0 ( .fault(fault), .net(N3883), .FEN(FEN[2260]), .op(N3883_t0) );
fim FAN_N3883_1 ( .fault(fault), .net(N3883), .FEN(FEN[2261]), .op(N3883_t1) );
fim FAN_N3889_0 ( .fault(fault), .net(N3889), .FEN(FEN[2262]), .op(N3889_t0) );
fim FAN_N3889_1 ( .fault(fault), .net(N3889), .FEN(FEN[2263]), .op(N3889_t1) );
fim FAN_N3889_2 ( .fault(fault), .net(N3889), .FEN(FEN[2264]), .op(N3889_t2) );
fim FAN_N3896_0 ( .fault(fault), .net(N3896), .FEN(FEN[2265]), .op(N3896_t0) );
fim FAN_N3896_1 ( .fault(fault), .net(N3896), .FEN(FEN[2266]), .op(N3896_t1) );
fim FAN_N3827_0 ( .fault(fault), .net(N3827), .FEN(FEN[2267]), .op(N3827_t0) );
fim FAN_N3827_1 ( .fault(fault), .net(N3827), .FEN(FEN[2268]), .op(N3827_t1) );
fim FAN_N3899_0 ( .fault(fault), .net(N3899), .FEN(FEN[2269]), .op(N3899_t0) );
fim FAN_N3899_1 ( .fault(fault), .net(N3899), .FEN(FEN[2270]), .op(N3899_t1) );
fim FAN_N3832_0 ( .fault(fault), .net(N3832), .FEN(FEN[2271]), .op(N3832_t0) );
fim FAN_N3832_1 ( .fault(fault), .net(N3832), .FEN(FEN[2272]), .op(N3832_t1) );
fim FAN_N3902_0 ( .fault(fault), .net(N3902), .FEN(FEN[2273]), .op(N3902_t0) );
fim FAN_N3902_1 ( .fault(fault), .net(N3902), .FEN(FEN[2274]), .op(N3902_t1) );
fim FAN_N3837_0 ( .fault(fault), .net(N3837), .FEN(FEN[2275]), .op(N3837_t0) );
fim FAN_N3837_1 ( .fault(fault), .net(N3837), .FEN(FEN[2276]), .op(N3837_t1) );
fim FAN_N3905_0 ( .fault(fault), .net(N3905), .FEN(FEN[2277]), .op(N3905_t0) );
fim FAN_N3905_1 ( .fault(fault), .net(N3905), .FEN(FEN[2278]), .op(N3905_t1) );
fim FAN_N3842_0 ( .fault(fault), .net(N3842), .FEN(FEN[2279]), .op(N3842_t0) );
fim FAN_N3842_1 ( .fault(fault), .net(N3842), .FEN(FEN[2280]), .op(N3842_t1) );
fim FAN_N3908_0 ( .fault(fault), .net(N3908), .FEN(FEN[2281]), .op(N3908_t0) );
fim FAN_N3908_1 ( .fault(fault), .net(N3908), .FEN(FEN[2282]), .op(N3908_t1) );
fim FAN_N3847_0 ( .fault(fault), .net(N3847), .FEN(FEN[2283]), .op(N3847_t0) );
fim FAN_N3847_1 ( .fault(fault), .net(N3847), .FEN(FEN[2284]), .op(N3847_t1) );
fim FAN_N3911_0 ( .fault(fault), .net(N3911), .FEN(FEN[2285]), .op(N3911_t0) );
fim FAN_N3911_1 ( .fault(fault), .net(N3911), .FEN(FEN[2286]), .op(N3911_t1) );
fim FAN_N3852_0 ( .fault(fault), .net(N3852), .FEN(FEN[2287]), .op(N3852_t0) );
fim FAN_N3852_1 ( .fault(fault), .net(N3852), .FEN(FEN[2288]), .op(N3852_t1) );
fim FAN_N3914_0 ( .fault(fault), .net(N3914), .FEN(FEN[2289]), .op(N3914_t0) );
fim FAN_N3914_1 ( .fault(fault), .net(N3914), .FEN(FEN[2290]), .op(N3914_t1) );
fim FAN_N3857_0 ( .fault(fault), .net(N3857), .FEN(FEN[2291]), .op(N3857_t0) );
fim FAN_N3857_1 ( .fault(fault), .net(N3857), .FEN(FEN[2292]), .op(N3857_t1) );
fim FAN_N3917_0 ( .fault(fault), .net(N3917), .FEN(FEN[2293]), .op(N3917_t0) );
fim FAN_N3917_1 ( .fault(fault), .net(N3917), .FEN(FEN[2294]), .op(N3917_t1) );
fim FAN_N3917_2 ( .fault(fault), .net(N3917), .FEN(FEN[2295]), .op(N3917_t2) );
fim FAN_N3923_0 ( .fault(fault), .net(N3923), .FEN(FEN[2296]), .op(N3923_t0) );
fim FAN_N3923_1 ( .fault(fault), .net(N3923), .FEN(FEN[2297]), .op(N3923_t1) );
fim FAN_N1002_0 ( .fault(fault), .net(N1002), .FEN(FEN[2298]), .op(N1002_t0) );
fim FAN_N1002_1 ( .fault(fault), .net(N1002), .FEN(FEN[2299]), .op(N1002_t1) );
fim FAN_N3926_0 ( .fault(fault), .net(N3926), .FEN(FEN[2300]), .op(N3926_t0) );
fim FAN_N3926_1 ( .fault(fault), .net(N3926), .FEN(FEN[2301]), .op(N3926_t1) );
fim FAN_N3926_2 ( .fault(fault), .net(N3926), .FEN(FEN[2302]), .op(N3926_t2) );
fim FAN_N3935_0 ( .fault(fault), .net(N3935), .FEN(FEN[2303]), .op(N3935_t0) );
fim FAN_N3935_1 ( .fault(fault), .net(N3935), .FEN(FEN[2304]), .op(N3935_t1) );
fim FAN_N3932_0 ( .fault(fault), .net(N3932), .FEN(FEN[2305]), .op(N3932_t0) );
fim FAN_N3932_1 ( .fault(fault), .net(N3932), .FEN(FEN[2306]), .op(N3932_t1) );
fim FAN_N3938_0 ( .fault(fault), .net(N3938), .FEN(FEN[2307]), .op(N3938_t0) );
fim FAN_N3938_1 ( .fault(fault), .net(N3938), .FEN(FEN[2308]), .op(N3938_t1) );
fim FAN_N3938_2 ( .fault(fault), .net(N3938), .FEN(FEN[2309]), .op(N3938_t2) );
fim FAN_N3944_0 ( .fault(fault), .net(N3944), .FEN(FEN[2310]), .op(N3944_t0) );
fim FAN_N3944_1 ( .fault(fault), .net(N3944), .FEN(FEN[2311]), .op(N3944_t1) );
fim FAN_N1245_0 ( .fault(fault), .net(N1245), .FEN(FEN[2312]), .op(N1245_t0) );
fim FAN_N1245_1 ( .fault(fault), .net(N1245), .FEN(FEN[2313]), .op(N1245_t1) );
fim FAN_N3947_0 ( .fault(fault), .net(N3947), .FEN(FEN[2314]), .op(N3947_t0) );
fim FAN_N3947_1 ( .fault(fault), .net(N3947), .FEN(FEN[2315]), .op(N3947_t1) );
fim FAN_N3947_2 ( .fault(fault), .net(N3947), .FEN(FEN[2316]), .op(N3947_t2) );
fim FAN_N3951_0 ( .fault(fault), .net(N3951), .FEN(FEN[2317]), .op(N3951_t0) );
fim FAN_N3951_1 ( .fault(fault), .net(N3951), .FEN(FEN[2318]), .op(N3951_t1) );
fim FAN_N3951_2 ( .fault(fault), .net(N3951), .FEN(FEN[2319]), .op(N3951_t2) );
fim FAN_N3955_0 ( .fault(fault), .net(N3955), .FEN(FEN[2320]), .op(N3955_t0) );
fim FAN_N3955_1 ( .fault(fault), .net(N3955), .FEN(FEN[2321]), .op(N3955_t1) );
fim FAN_N3955_2 ( .fault(fault), .net(N3955), .FEN(FEN[2322]), .op(N3955_t2) );
fim FAN_N3959_0 ( .fault(fault), .net(N3959), .FEN(FEN[2323]), .op(N3959_t0) );
fim FAN_N3959_1 ( .fault(fault), .net(N3959), .FEN(FEN[2324]), .op(N3959_t1) );
fim FAN_N3959_2 ( .fault(fault), .net(N3959), .FEN(FEN[2325]), .op(N3959_t2) );
fim FAN_N3963_0 ( .fault(fault), .net(N3963), .FEN(FEN[2326]), .op(N3963_t0) );
fim FAN_N3963_1 ( .fault(fault), .net(N3963), .FEN(FEN[2327]), .op(N3963_t1) );
fim FAN_N3963_2 ( .fault(fault), .net(N3963), .FEN(FEN[2328]), .op(N3963_t2) );
fim FAN_N3967_0 ( .fault(fault), .net(N3967), .FEN(FEN[2329]), .op(N3967_t0) );
fim FAN_N3967_1 ( .fault(fault), .net(N3967), .FEN(FEN[2330]), .op(N3967_t1) );
fim FAN_N3967_2 ( .fault(fault), .net(N3967), .FEN(FEN[2331]), .op(N3967_t2) );
fim FAN_N3971_0 ( .fault(fault), .net(N3971), .FEN(FEN[2332]), .op(N3971_t0) );
fim FAN_N3971_1 ( .fault(fault), .net(N3971), .FEN(FEN[2333]), .op(N3971_t1) );
fim FAN_N3971_2 ( .fault(fault), .net(N3971), .FEN(FEN[2334]), .op(N3971_t2) );
fim FAN_N3977_0 ( .fault(fault), .net(N3977), .FEN(FEN[2335]), .op(N3977_t0) );
fim FAN_N3977_1 ( .fault(fault), .net(N3977), .FEN(FEN[2336]), .op(N3977_t1) );
fim FAN_N954_0 ( .fault(fault), .net(N954), .FEN(FEN[2337]), .op(N954_t0) );
fim FAN_N954_1 ( .fault(fault), .net(N954), .FEN(FEN[2338]), .op(N954_t1) );
fim FAN_N3980_0 ( .fault(fault), .net(N3980), .FEN(FEN[2339]), .op(N3980_t0) );
fim FAN_N3980_1 ( .fault(fault), .net(N3980), .FEN(FEN[2340]), .op(N3980_t1) );
fim FAN_N3980_2 ( .fault(fault), .net(N3980), .FEN(FEN[2341]), .op(N3980_t2) );
fim FAN_N3989_0 ( .fault(fault), .net(N3989), .FEN(FEN[2342]), .op(N3989_t0) );
fim FAN_N3989_1 ( .fault(fault), .net(N3989), .FEN(FEN[2343]), .op(N3989_t1) );
fim FAN_N3986_0 ( .fault(fault), .net(N3986), .FEN(FEN[2344]), .op(N3986_t0) );
fim FAN_N3986_1 ( .fault(fault), .net(N3986), .FEN(FEN[2345]), .op(N3986_t1) );
fim FAN_N3992_0 ( .fault(fault), .net(N3992), .FEN(FEN[2346]), .op(N3992_t0) );
fim FAN_N3992_1 ( .fault(fault), .net(N3992), .FEN(FEN[2347]), .op(N3992_t1) );
fim FAN_N3992_2 ( .fault(fault), .net(N3992), .FEN(FEN[2348]), .op(N3992_t2) );
fim FAN_N3998_0 ( .fault(fault), .net(N3998), .FEN(FEN[2349]), .op(N3998_t0) );
fim FAN_N3998_1 ( .fault(fault), .net(N3998), .FEN(FEN[2350]), .op(N3998_t1) );
fim FAN_N1197_0 ( .fault(fault), .net(N1197), .FEN(FEN[2351]), .op(N1197_t0) );
fim FAN_N1197_1 ( .fault(fault), .net(N1197), .FEN(FEN[2352]), .op(N1197_t1) );
fim FAN_N4001_0 ( .fault(fault), .net(N4001), .FEN(FEN[2353]), .op(N4001_t0) );
fim FAN_N4001_1 ( .fault(fault), .net(N4001), .FEN(FEN[2354]), .op(N4001_t1) );
fim FAN_N4001_2 ( .fault(fault), .net(N4001), .FEN(FEN[2355]), .op(N4001_t2) );
fim FAN_N4019_0 ( .fault(fault), .net(N4019), .FEN(FEN[2356]), .op(N4019_t0) );
fim FAN_N4019_1 ( .fault(fault), .net(N4019), .FEN(FEN[2357]), .op(N4019_t1) );
fim FAN_N906_0 ( .fault(fault), .net(N906), .FEN(FEN[2358]), .op(N906_t0) );
fim FAN_N906_1 ( .fault(fault), .net(N906), .FEN(FEN[2359]), .op(N906_t1) );
fim FAN_N4022_0 ( .fault(fault), .net(N4022), .FEN(FEN[2360]), .op(N4022_t0) );
fim FAN_N4022_1 ( .fault(fault), .net(N4022), .FEN(FEN[2361]), .op(N4022_t1) );
fim FAN_N4022_2 ( .fault(fault), .net(N4022), .FEN(FEN[2362]), .op(N4022_t2) );
fim FAN_N4031_0 ( .fault(fault), .net(N4031), .FEN(FEN[2363]), .op(N4031_t0) );
fim FAN_N4031_1 ( .fault(fault), .net(N4031), .FEN(FEN[2364]), .op(N4031_t1) );
fim FAN_N4028_0 ( .fault(fault), .net(N4028), .FEN(FEN[2365]), .op(N4028_t0) );
fim FAN_N4028_1 ( .fault(fault), .net(N4028), .FEN(FEN[2366]), .op(N4028_t1) );
fim FAN_N4034_0 ( .fault(fault), .net(N4034), .FEN(FEN[2367]), .op(N4034_t0) );
fim FAN_N4034_1 ( .fault(fault), .net(N4034), .FEN(FEN[2368]), .op(N4034_t1) );
fim FAN_N4034_2 ( .fault(fault), .net(N4034), .FEN(FEN[2369]), .op(N4034_t2) );
fim FAN_N4040_0 ( .fault(fault), .net(N4040), .FEN(FEN[2370]), .op(N4040_t0) );
fim FAN_N4040_1 ( .fault(fault), .net(N4040), .FEN(FEN[2371]), .op(N4040_t1) );
fim FAN_N1149_0 ( .fault(fault), .net(N1149), .FEN(FEN[2372]), .op(N1149_t0) );
fim FAN_N1149_1 ( .fault(fault), .net(N1149), .FEN(FEN[2373]), .op(N1149_t1) );
fim FAN_N4043_0 ( .fault(fault), .net(N4043), .FEN(FEN[2374]), .op(N4043_t0) );
fim FAN_N4043_1 ( .fault(fault), .net(N4043), .FEN(FEN[2375]), .op(N4043_t1) );
fim FAN_N4043_2 ( .fault(fault), .net(N4043), .FEN(FEN[2376]), .op(N4043_t2) );
fim FAN_N1293_0 ( .fault(fault), .net(N1293), .FEN(FEN[2377]), .op(N1293_t0) );
fim FAN_N1293_1 ( .fault(fault), .net(N1293), .FEN(FEN[2378]), .op(N1293_t1) );
fim FAN_N4049_0 ( .fault(fault), .net(N4049), .FEN(FEN[2379]), .op(N4049_t0) );
fim FAN_N4049_1 ( .fault(fault), .net(N4049), .FEN(FEN[2380]), .op(N4049_t1) );
fim FAN_N4052_0 ( .fault(fault), .net(N4052), .FEN(FEN[2381]), .op(N4052_t0) );
fim FAN_N4052_1 ( .fault(fault), .net(N4052), .FEN(FEN[2382]), .op(N4052_t1) );
fim FAN_N570_0 ( .fault(fault), .net(N570), .FEN(FEN[2383]), .op(N570_t0) );
fim FAN_N570_1 ( .fault(fault), .net(N570), .FEN(FEN[2384]), .op(N570_t1) );
fim FAN_N4055_0 ( .fault(fault), .net(N4055), .FEN(FEN[2385]), .op(N4055_t0) );
fim FAN_N4055_1 ( .fault(fault), .net(N4055), .FEN(FEN[2386]), .op(N4055_t1) );
fim FAN_N618_0 ( .fault(fault), .net(N618), .FEN(FEN[2387]), .op(N618_t0) );
fim FAN_N618_1 ( .fault(fault), .net(N618), .FEN(FEN[2388]), .op(N618_t1) );
fim FAN_N4058_0 ( .fault(fault), .net(N4058), .FEN(FEN[2389]), .op(N4058_t0) );
fim FAN_N4058_1 ( .fault(fault), .net(N4058), .FEN(FEN[2390]), .op(N4058_t1) );
fim FAN_N666_0 ( .fault(fault), .net(N666), .FEN(FEN[2391]), .op(N666_t0) );
fim FAN_N666_1 ( .fault(fault), .net(N666), .FEN(FEN[2392]), .op(N666_t1) );
fim FAN_N4061_0 ( .fault(fault), .net(N4061), .FEN(FEN[2393]), .op(N4061_t0) );
fim FAN_N4061_1 ( .fault(fault), .net(N4061), .FEN(FEN[2394]), .op(N4061_t1) );
fim FAN_N714_0 ( .fault(fault), .net(N714), .FEN(FEN[2395]), .op(N714_t0) );
fim FAN_N714_1 ( .fault(fault), .net(N714), .FEN(FEN[2396]), .op(N714_t1) );
fim FAN_N4064_0 ( .fault(fault), .net(N4064), .FEN(FEN[2397]), .op(N4064_t0) );
fim FAN_N4064_1 ( .fault(fault), .net(N4064), .FEN(FEN[2398]), .op(N4064_t1) );
fim FAN_N762_0 ( .fault(fault), .net(N762), .FEN(FEN[2399]), .op(N762_t0) );
fim FAN_N762_1 ( .fault(fault), .net(N762), .FEN(FEN[2400]), .op(N762_t1) );
fim FAN_N4067_0 ( .fault(fault), .net(N4067), .FEN(FEN[2401]), .op(N4067_t0) );
fim FAN_N4067_1 ( .fault(fault), .net(N4067), .FEN(FEN[2402]), .op(N4067_t1) );
fim FAN_N810_0 ( .fault(fault), .net(N810), .FEN(FEN[2403]), .op(N810_t0) );
fim FAN_N810_1 ( .fault(fault), .net(N810), .FEN(FEN[2404]), .op(N810_t1) );
fim FAN_N4070_0 ( .fault(fault), .net(N4070), .FEN(FEN[2405]), .op(N4070_t0) );
fim FAN_N4070_1 ( .fault(fault), .net(N4070), .FEN(FEN[2406]), .op(N4070_t1) );
fim FAN_N858_0 ( .fault(fault), .net(N858), .FEN(FEN[2407]), .op(N858_t0) );
fim FAN_N858_1 ( .fault(fault), .net(N858), .FEN(FEN[2408]), .op(N858_t1) );
fim FAN_N4073_0 ( .fault(fault), .net(N4073), .FEN(FEN[2409]), .op(N4073_t0) );
fim FAN_N4073_1 ( .fault(fault), .net(N4073), .FEN(FEN[2410]), .op(N4073_t1) );
fim FAN_N4073_2 ( .fault(fault), .net(N4073), .FEN(FEN[2411]), .op(N4073_t2) );
fim FAN_N4082_0 ( .fault(fault), .net(N4082), .FEN(FEN[2412]), .op(N4082_t0) );
fim FAN_N4082_1 ( .fault(fault), .net(N4082), .FEN(FEN[2413]), .op(N4082_t1) );
fim FAN_N4079_0 ( .fault(fault), .net(N4079), .FEN(FEN[2414]), .op(N4079_t0) );
fim FAN_N4079_1 ( .fault(fault), .net(N4079), .FEN(FEN[2415]), .op(N4079_t1) );
fim FAN_N4085_0 ( .fault(fault), .net(N4085), .FEN(FEN[2416]), .op(N4085_t0) );
fim FAN_N4085_1 ( .fault(fault), .net(N4085), .FEN(FEN[2417]), .op(N4085_t1) );
fim FAN_N4085_2 ( .fault(fault), .net(N4085), .FEN(FEN[2418]), .op(N4085_t2) );
fim FAN_N4091_0 ( .fault(fault), .net(N4091), .FEN(FEN[2419]), .op(N4091_t0) );
fim FAN_N4091_1 ( .fault(fault), .net(N4091), .FEN(FEN[2420]), .op(N4091_t1) );
fim FAN_N1101_0 ( .fault(fault), .net(N1101), .FEN(FEN[2421]), .op(N1101_t0) );
fim FAN_N1101_1 ( .fault(fault), .net(N1101), .FEN(FEN[2422]), .op(N1101_t1) );
fim FAN_N4094_0 ( .fault(fault), .net(N4094), .FEN(FEN[2423]), .op(N4094_t0) );
fim FAN_N4094_1 ( .fault(fault), .net(N4094), .FEN(FEN[2424]), .op(N4094_t1) );
fim FAN_N4094_2 ( .fault(fault), .net(N4094), .FEN(FEN[2425]), .op(N4094_t2) );
fim FAN_N4103_0 ( .fault(fault), .net(N4103), .FEN(FEN[2426]), .op(N4103_t0) );
fim FAN_N4103_1 ( .fault(fault), .net(N4103), .FEN(FEN[2427]), .op(N4103_t1) );
fim FAN_N4100_0 ( .fault(fault), .net(N4100), .FEN(FEN[2428]), .op(N4100_t0) );
fim FAN_N4100_1 ( .fault(fault), .net(N4100), .FEN(FEN[2429]), .op(N4100_t1) );
fim FAN_N4106_0 ( .fault(fault), .net(N4106), .FEN(FEN[2430]), .op(N4106_t0) );
fim FAN_N4106_1 ( .fault(fault), .net(N4106), .FEN(FEN[2431]), .op(N4106_t1) );
fim FAN_N4106_2 ( .fault(fault), .net(N4106), .FEN(FEN[2432]), .op(N4106_t2) );
fim FAN_N4110_0 ( .fault(fault), .net(N4110), .FEN(FEN[2433]), .op(N4110_t0) );
fim FAN_N4110_1 ( .fault(fault), .net(N4110), .FEN(FEN[2434]), .op(N4110_t1) );
fim FAN_N4110_2 ( .fault(fault), .net(N4110), .FEN(FEN[2435]), .op(N4110_t2) );
fim FAN_N4114_0 ( .fault(fault), .net(N4114), .FEN(FEN[2436]), .op(N4114_t0) );
fim FAN_N4114_1 ( .fault(fault), .net(N4114), .FEN(FEN[2437]), .op(N4114_t1) );
fim FAN_N4114_2 ( .fault(fault), .net(N4114), .FEN(FEN[2438]), .op(N4114_t2) );
fim FAN_N4118_0 ( .fault(fault), .net(N4118), .FEN(FEN[2439]), .op(N4118_t0) );
fim FAN_N4118_1 ( .fault(fault), .net(N4118), .FEN(FEN[2440]), .op(N4118_t1) );
fim FAN_N4118_2 ( .fault(fault), .net(N4118), .FEN(FEN[2441]), .op(N4118_t2) );
fim FAN_N4122_0 ( .fault(fault), .net(N4122), .FEN(FEN[2442]), .op(N4122_t0) );
fim FAN_N4122_1 ( .fault(fault), .net(N4122), .FEN(FEN[2443]), .op(N4122_t1) );
fim FAN_N4122_2 ( .fault(fault), .net(N4122), .FEN(FEN[2444]), .op(N4122_t2) );
fim FAN_N4126_0 ( .fault(fault), .net(N4126), .FEN(FEN[2445]), .op(N4126_t0) );
fim FAN_N4126_1 ( .fault(fault), .net(N4126), .FEN(FEN[2446]), .op(N4126_t1) );
fim FAN_N4126_2 ( .fault(fault), .net(N4126), .FEN(FEN[2447]), .op(N4126_t2) );
fim FAN_N4130_0 ( .fault(fault), .net(N4130), .FEN(FEN[2448]), .op(N4130_t0) );
fim FAN_N4130_1 ( .fault(fault), .net(N4130), .FEN(FEN[2449]), .op(N4130_t1) );
fim FAN_N4130_2 ( .fault(fault), .net(N4130), .FEN(FEN[2450]), .op(N4130_t2) );
fim FAN_N4134_0 ( .fault(fault), .net(N4134), .FEN(FEN[2451]), .op(N4134_t0) );
fim FAN_N4134_1 ( .fault(fault), .net(N4134), .FEN(FEN[2452]), .op(N4134_t1) );
fim FAN_N4134_2 ( .fault(fault), .net(N4134), .FEN(FEN[2453]), .op(N4134_t2) );
fim FAN_N4143_0 ( .fault(fault), .net(N4143), .FEN(FEN[2454]), .op(N4143_t0) );
fim FAN_N4143_1 ( .fault(fault), .net(N4143), .FEN(FEN[2455]), .op(N4143_t1) );
fim FAN_N4140_0 ( .fault(fault), .net(N4140), .FEN(FEN[2456]), .op(N4140_t0) );
fim FAN_N4140_1 ( .fault(fault), .net(N4140), .FEN(FEN[2457]), .op(N4140_t1) );
fim FAN_N4146_0 ( .fault(fault), .net(N4146), .FEN(FEN[2458]), .op(N4146_t0) );
fim FAN_N4146_1 ( .fault(fault), .net(N4146), .FEN(FEN[2459]), .op(N4146_t1) );
fim FAN_N4146_2 ( .fault(fault), .net(N4146), .FEN(FEN[2460]), .op(N4146_t2) );
fim FAN_N4152_0 ( .fault(fault), .net(N4152), .FEN(FEN[2461]), .op(N4152_t0) );
fim FAN_N4152_1 ( .fault(fault), .net(N4152), .FEN(FEN[2462]), .op(N4152_t1) );
fim FAN_N1053_0 ( .fault(fault), .net(N1053), .FEN(FEN[2463]), .op(N1053_t0) );
fim FAN_N1053_1 ( .fault(fault), .net(N1053), .FEN(FEN[2464]), .op(N1053_t1) );
fim FAN_N4155_0 ( .fault(fault), .net(N4155), .FEN(FEN[2465]), .op(N4155_t0) );
fim FAN_N4155_1 ( .fault(fault), .net(N4155), .FEN(FEN[2466]), .op(N4155_t1) );
fim FAN_N4155_2 ( .fault(fault), .net(N4155), .FEN(FEN[2467]), .op(N4155_t2) );
fim FAN_N4164_0 ( .fault(fault), .net(N4164), .FEN(FEN[2468]), .op(N4164_t0) );
fim FAN_N4164_1 ( .fault(fault), .net(N4164), .FEN(FEN[2469]), .op(N4164_t1) );
fim FAN_N4161_0 ( .fault(fault), .net(N4161), .FEN(FEN[2470]), .op(N4161_t0) );
fim FAN_N4161_1 ( .fault(fault), .net(N4161), .FEN(FEN[2471]), .op(N4161_t1) );
fim FAN_N4167_0 ( .fault(fault), .net(N4167), .FEN(FEN[2472]), .op(N4167_t0) );
fim FAN_N4167_1 ( .fault(fault), .net(N4167), .FEN(FEN[2473]), .op(N4167_t1) );
fim FAN_N4167_2 ( .fault(fault), .net(N4167), .FEN(FEN[2474]), .op(N4167_t2) );
fim FAN_N4208_0 ( .fault(fault), .net(N4208), .FEN(FEN[2475]), .op(N4208_t0) );
fim FAN_N4208_1 ( .fault(fault), .net(N4208), .FEN(FEN[2476]), .op(N4208_t1) );
fim FAN_N4205_0 ( .fault(fault), .net(N4205), .FEN(FEN[2477]), .op(N4205_t0) );
fim FAN_N4205_1 ( .fault(fault), .net(N4205), .FEN(FEN[2478]), .op(N4205_t1) );
fim FAN_N4211_0 ( .fault(fault), .net(N4211), .FEN(FEN[2479]), .op(N4211_t0) );
fim FAN_N4211_1 ( .fault(fault), .net(N4211), .FEN(FEN[2480]), .op(N4211_t1) );
fim FAN_N4211_2 ( .fault(fault), .net(N4211), .FEN(FEN[2481]), .op(N4211_t2) );
fim FAN_N4217_0 ( .fault(fault), .net(N4217), .FEN(FEN[2482]), .op(N4217_t0) );
fim FAN_N4217_1 ( .fault(fault), .net(N4217), .FEN(FEN[2483]), .op(N4217_t1) );
fim FAN_N1005_0 ( .fault(fault), .net(N1005), .FEN(FEN[2484]), .op(N1005_t0) );
fim FAN_N1005_1 ( .fault(fault), .net(N1005), .FEN(FEN[2485]), .op(N1005_t1) );
fim FAN_N4220_0 ( .fault(fault), .net(N4220), .FEN(FEN[2486]), .op(N4220_t0) );
fim FAN_N4220_1 ( .fault(fault), .net(N4220), .FEN(FEN[2487]), .op(N4220_t1) );
fim FAN_N4220_2 ( .fault(fault), .net(N4220), .FEN(FEN[2488]), .op(N4220_t2) );
fim FAN_N4229_0 ( .fault(fault), .net(N4229), .FEN(FEN[2489]), .op(N4229_t0) );
fim FAN_N4229_1 ( .fault(fault), .net(N4229), .FEN(FEN[2490]), .op(N4229_t1) );
fim FAN_N4226_0 ( .fault(fault), .net(N4226), .FEN(FEN[2491]), .op(N4226_t0) );
fim FAN_N4226_1 ( .fault(fault), .net(N4226), .FEN(FEN[2492]), .op(N4226_t1) );
fim FAN_N4232_0 ( .fault(fault), .net(N4232), .FEN(FEN[2493]), .op(N4232_t0) );
fim FAN_N4232_1 ( .fault(fault), .net(N4232), .FEN(FEN[2494]), .op(N4232_t1) );
fim FAN_N4232_2 ( .fault(fault), .net(N4232), .FEN(FEN[2495]), .op(N4232_t2) );
fim FAN_N4238_0 ( .fault(fault), .net(N4238), .FEN(FEN[2496]), .op(N4238_t0) );
fim FAN_N4238_1 ( .fault(fault), .net(N4238), .FEN(FEN[2497]), .op(N4238_t1) );
fim FAN_N1248_0 ( .fault(fault), .net(N1248), .FEN(FEN[2498]), .op(N1248_t0) );
fim FAN_N1248_1 ( .fault(fault), .net(N1248), .FEN(FEN[2499]), .op(N1248_t1) );
fim FAN_N4242_0 ( .fault(fault), .net(N4242), .FEN(FEN[2500]), .op(N4242_t0) );
fim FAN_N4242_1 ( .fault(fault), .net(N4242), .FEN(FEN[2501]), .op(N4242_t1) );
fim FAN_N4175_0 ( .fault(fault), .net(N4175), .FEN(FEN[2502]), .op(N4175_t0) );
fim FAN_N4175_1 ( .fault(fault), .net(N4175), .FEN(FEN[2503]), .op(N4175_t1) );
fim FAN_N4245_0 ( .fault(fault), .net(N4245), .FEN(FEN[2504]), .op(N4245_t0) );
fim FAN_N4245_1 ( .fault(fault), .net(N4245), .FEN(FEN[2505]), .op(N4245_t1) );
fim FAN_N4180_0 ( .fault(fault), .net(N4180), .FEN(FEN[2506]), .op(N4180_t0) );
fim FAN_N4180_1 ( .fault(fault), .net(N4180), .FEN(FEN[2507]), .op(N4180_t1) );
fim FAN_N4248_0 ( .fault(fault), .net(N4248), .FEN(FEN[2508]), .op(N4248_t0) );
fim FAN_N4248_1 ( .fault(fault), .net(N4248), .FEN(FEN[2509]), .op(N4248_t1) );
fim FAN_N4185_0 ( .fault(fault), .net(N4185), .FEN(FEN[2510]), .op(N4185_t0) );
fim FAN_N4185_1 ( .fault(fault), .net(N4185), .FEN(FEN[2511]), .op(N4185_t1) );
fim FAN_N4251_0 ( .fault(fault), .net(N4251), .FEN(FEN[2512]), .op(N4251_t0) );
fim FAN_N4251_1 ( .fault(fault), .net(N4251), .FEN(FEN[2513]), .op(N4251_t1) );
fim FAN_N4190_0 ( .fault(fault), .net(N4190), .FEN(FEN[2514]), .op(N4190_t0) );
fim FAN_N4190_1 ( .fault(fault), .net(N4190), .FEN(FEN[2515]), .op(N4190_t1) );
fim FAN_N4254_0 ( .fault(fault), .net(N4254), .FEN(FEN[2516]), .op(N4254_t0) );
fim FAN_N4254_1 ( .fault(fault), .net(N4254), .FEN(FEN[2517]), .op(N4254_t1) );
fim FAN_N4195_0 ( .fault(fault), .net(N4195), .FEN(FEN[2518]), .op(N4195_t0) );
fim FAN_N4195_1 ( .fault(fault), .net(N4195), .FEN(FEN[2519]), .op(N4195_t1) );
fim FAN_N4257_0 ( .fault(fault), .net(N4257), .FEN(FEN[2520]), .op(N4257_t0) );
fim FAN_N4257_1 ( .fault(fault), .net(N4257), .FEN(FEN[2521]), .op(N4257_t1) );
fim FAN_N4200_0 ( .fault(fault), .net(N4200), .FEN(FEN[2522]), .op(N4200_t0) );
fim FAN_N4200_1 ( .fault(fault), .net(N4200), .FEN(FEN[2523]), .op(N4200_t1) );
fim FAN_N4260_0 ( .fault(fault), .net(N4260), .FEN(FEN[2524]), .op(N4260_t0) );
fim FAN_N4260_1 ( .fault(fault), .net(N4260), .FEN(FEN[2525]), .op(N4260_t1) );
fim FAN_N4260_2 ( .fault(fault), .net(N4260), .FEN(FEN[2526]), .op(N4260_t2) );
fim FAN_N4266_0 ( .fault(fault), .net(N4266), .FEN(FEN[2527]), .op(N4266_t0) );
fim FAN_N4266_1 ( .fault(fault), .net(N4266), .FEN(FEN[2528]), .op(N4266_t1) );
fim FAN_N957_0 ( .fault(fault), .net(N957), .FEN(FEN[2529]), .op(N957_t0) );
fim FAN_N957_1 ( .fault(fault), .net(N957), .FEN(FEN[2530]), .op(N957_t1) );
fim FAN_N4269_0 ( .fault(fault), .net(N4269), .FEN(FEN[2531]), .op(N4269_t0) );
fim FAN_N4269_1 ( .fault(fault), .net(N4269), .FEN(FEN[2532]), .op(N4269_t1) );
fim FAN_N4269_2 ( .fault(fault), .net(N4269), .FEN(FEN[2533]), .op(N4269_t2) );
fim FAN_N4278_0 ( .fault(fault), .net(N4278), .FEN(FEN[2534]), .op(N4278_t0) );
fim FAN_N4278_1 ( .fault(fault), .net(N4278), .FEN(FEN[2535]), .op(N4278_t1) );
fim FAN_N4275_0 ( .fault(fault), .net(N4275), .FEN(FEN[2536]), .op(N4275_t0) );
fim FAN_N4275_1 ( .fault(fault), .net(N4275), .FEN(FEN[2537]), .op(N4275_t1) );
fim FAN_N4281_0 ( .fault(fault), .net(N4281), .FEN(FEN[2538]), .op(N4281_t0) );
fim FAN_N4281_1 ( .fault(fault), .net(N4281), .FEN(FEN[2539]), .op(N4281_t1) );
fim FAN_N4281_2 ( .fault(fault), .net(N4281), .FEN(FEN[2540]), .op(N4281_t2) );
fim FAN_N4287_0 ( .fault(fault), .net(N4287), .FEN(FEN[2541]), .op(N4287_t0) );
fim FAN_N4287_1 ( .fault(fault), .net(N4287), .FEN(FEN[2542]), .op(N4287_t1) );
fim FAN_N1200_0 ( .fault(fault), .net(N1200), .FEN(FEN[2543]), .op(N1200_t0) );
fim FAN_N1200_1 ( .fault(fault), .net(N1200), .FEN(FEN[2544]), .op(N1200_t1) );
fim FAN_N4290_0 ( .fault(fault), .net(N4290), .FEN(FEN[2545]), .op(N4290_t0) );
fim FAN_N4290_1 ( .fault(fault), .net(N4290), .FEN(FEN[2546]), .op(N4290_t1) );
fim FAN_N4290_2 ( .fault(fault), .net(N4290), .FEN(FEN[2547]), .op(N4290_t2) );
fim FAN_N4294_0 ( .fault(fault), .net(N4294), .FEN(FEN[2548]), .op(N4294_t0) );
fim FAN_N4294_1 ( .fault(fault), .net(N4294), .FEN(FEN[2549]), .op(N4294_t1) );
fim FAN_N4294_2 ( .fault(fault), .net(N4294), .FEN(FEN[2550]), .op(N4294_t2) );
fim FAN_N4298_0 ( .fault(fault), .net(N4298), .FEN(FEN[2551]), .op(N4298_t0) );
fim FAN_N4298_1 ( .fault(fault), .net(N4298), .FEN(FEN[2552]), .op(N4298_t1) );
fim FAN_N4298_2 ( .fault(fault), .net(N4298), .FEN(FEN[2553]), .op(N4298_t2) );
fim FAN_N4302_0 ( .fault(fault), .net(N4302), .FEN(FEN[2554]), .op(N4302_t0) );
fim FAN_N4302_1 ( .fault(fault), .net(N4302), .FEN(FEN[2555]), .op(N4302_t1) );
fim FAN_N4302_2 ( .fault(fault), .net(N4302), .FEN(FEN[2556]), .op(N4302_t2) );
fim FAN_N4306_0 ( .fault(fault), .net(N4306), .FEN(FEN[2557]), .op(N4306_t0) );
fim FAN_N4306_1 ( .fault(fault), .net(N4306), .FEN(FEN[2558]), .op(N4306_t1) );
fim FAN_N4306_2 ( .fault(fault), .net(N4306), .FEN(FEN[2559]), .op(N4306_t2) );
fim FAN_N4310_0 ( .fault(fault), .net(N4310), .FEN(FEN[2560]), .op(N4310_t0) );
fim FAN_N4310_1 ( .fault(fault), .net(N4310), .FEN(FEN[2561]), .op(N4310_t1) );
fim FAN_N4310_2 ( .fault(fault), .net(N4310), .FEN(FEN[2562]), .op(N4310_t2) );
fim FAN_N4314_0 ( .fault(fault), .net(N4314), .FEN(FEN[2563]), .op(N4314_t0) );
fim FAN_N4314_1 ( .fault(fault), .net(N4314), .FEN(FEN[2564]), .op(N4314_t1) );
fim FAN_N4314_2 ( .fault(fault), .net(N4314), .FEN(FEN[2565]), .op(N4314_t2) );
fim FAN_N4320_0 ( .fault(fault), .net(N4320), .FEN(FEN[2566]), .op(N4320_t0) );
fim FAN_N4320_1 ( .fault(fault), .net(N4320), .FEN(FEN[2567]), .op(N4320_t1) );
fim FAN_N909_0 ( .fault(fault), .net(N909), .FEN(FEN[2568]), .op(N909_t0) );
fim FAN_N909_1 ( .fault(fault), .net(N909), .FEN(FEN[2569]), .op(N909_t1) );
fim FAN_N4323_0 ( .fault(fault), .net(N4323), .FEN(FEN[2570]), .op(N4323_t0) );
fim FAN_N4323_1 ( .fault(fault), .net(N4323), .FEN(FEN[2571]), .op(N4323_t1) );
fim FAN_N4323_2 ( .fault(fault), .net(N4323), .FEN(FEN[2572]), .op(N4323_t2) );
fim FAN_N4332_0 ( .fault(fault), .net(N4332), .FEN(FEN[2573]), .op(N4332_t0) );
fim FAN_N4332_1 ( .fault(fault), .net(N4332), .FEN(FEN[2574]), .op(N4332_t1) );
fim FAN_N4329_0 ( .fault(fault), .net(N4329), .FEN(FEN[2575]), .op(N4329_t0) );
fim FAN_N4329_1 ( .fault(fault), .net(N4329), .FEN(FEN[2576]), .op(N4329_t1) );
fim FAN_N4335_0 ( .fault(fault), .net(N4335), .FEN(FEN[2577]), .op(N4335_t0) );
fim FAN_N4335_1 ( .fault(fault), .net(N4335), .FEN(FEN[2578]), .op(N4335_t1) );
fim FAN_N4335_2 ( .fault(fault), .net(N4335), .FEN(FEN[2579]), .op(N4335_t2) );
fim FAN_N4341_0 ( .fault(fault), .net(N4341), .FEN(FEN[2580]), .op(N4341_t0) );
fim FAN_N4341_1 ( .fault(fault), .net(N4341), .FEN(FEN[2581]), .op(N4341_t1) );
fim FAN_N1152_0 ( .fault(fault), .net(N1152), .FEN(FEN[2582]), .op(N1152_t0) );
fim FAN_N1152_1 ( .fault(fault), .net(N1152), .FEN(FEN[2583]), .op(N1152_t1) );
fim FAN_N4344_0 ( .fault(fault), .net(N4344), .FEN(FEN[2584]), .op(N4344_t0) );
fim FAN_N4344_1 ( .fault(fault), .net(N4344), .FEN(FEN[2585]), .op(N4344_t1) );
fim FAN_N4344_2 ( .fault(fault), .net(N4344), .FEN(FEN[2586]), .op(N4344_t2) );
fim FAN_N1296_0 ( .fault(fault), .net(N1296), .FEN(FEN[2587]), .op(N1296_t0) );
fim FAN_N1296_1 ( .fault(fault), .net(N1296), .FEN(FEN[2588]), .op(N1296_t1) );
fim FAN_N4350_0 ( .fault(fault), .net(N4350), .FEN(FEN[2589]), .op(N4350_t0) );
fim FAN_N4350_1 ( .fault(fault), .net(N4350), .FEN(FEN[2590]), .op(N4350_t1) );
fim FAN_N4365_0 ( .fault(fault), .net(N4365), .FEN(FEN[2591]), .op(N4365_t0) );
fim FAN_N4365_1 ( .fault(fault), .net(N4365), .FEN(FEN[2592]), .op(N4365_t1) );
fim FAN_N861_0 ( .fault(fault), .net(N861), .FEN(FEN[2593]), .op(N861_t0) );
fim FAN_N861_1 ( .fault(fault), .net(N861), .FEN(FEN[2594]), .op(N861_t1) );
fim FAN_N4368_0 ( .fault(fault), .net(N4368), .FEN(FEN[2595]), .op(N4368_t0) );
fim FAN_N4368_1 ( .fault(fault), .net(N4368), .FEN(FEN[2596]), .op(N4368_t1) );
fim FAN_N4368_2 ( .fault(fault), .net(N4368), .FEN(FEN[2597]), .op(N4368_t2) );
fim FAN_N4377_0 ( .fault(fault), .net(N4377), .FEN(FEN[2598]), .op(N4377_t0) );
fim FAN_N4377_1 ( .fault(fault), .net(N4377), .FEN(FEN[2599]), .op(N4377_t1) );
fim FAN_N4374_0 ( .fault(fault), .net(N4374), .FEN(FEN[2600]), .op(N4374_t0) );
fim FAN_N4374_1 ( .fault(fault), .net(N4374), .FEN(FEN[2601]), .op(N4374_t1) );
fim FAN_N4380_0 ( .fault(fault), .net(N4380), .FEN(FEN[2602]), .op(N4380_t0) );
fim FAN_N4380_1 ( .fault(fault), .net(N4380), .FEN(FEN[2603]), .op(N4380_t1) );
fim FAN_N4380_2 ( .fault(fault), .net(N4380), .FEN(FEN[2604]), .op(N4380_t2) );
fim FAN_N4386_0 ( .fault(fault), .net(N4386), .FEN(FEN[2605]), .op(N4386_t0) );
fim FAN_N4386_1 ( .fault(fault), .net(N4386), .FEN(FEN[2606]), .op(N4386_t1) );
fim FAN_N1104_0 ( .fault(fault), .net(N1104), .FEN(FEN[2607]), .op(N1104_t0) );
fim FAN_N1104_1 ( .fault(fault), .net(N1104), .FEN(FEN[2608]), .op(N1104_t1) );
fim FAN_N4389_0 ( .fault(fault), .net(N4389), .FEN(FEN[2609]), .op(N4389_t0) );
fim FAN_N4389_1 ( .fault(fault), .net(N4389), .FEN(FEN[2610]), .op(N4389_t1) );
fim FAN_N4389_2 ( .fault(fault), .net(N4389), .FEN(FEN[2611]), .op(N4389_t2) );
fim FAN_N4398_0 ( .fault(fault), .net(N4398), .FEN(FEN[2612]), .op(N4398_t0) );
fim FAN_N4398_1 ( .fault(fault), .net(N4398), .FEN(FEN[2613]), .op(N4398_t1) );
fim FAN_N4395_0 ( .fault(fault), .net(N4395), .FEN(FEN[2614]), .op(N4395_t0) );
fim FAN_N4395_1 ( .fault(fault), .net(N4395), .FEN(FEN[2615]), .op(N4395_t1) );
fim FAN_N4401_0 ( .fault(fault), .net(N4401), .FEN(FEN[2616]), .op(N4401_t0) );
fim FAN_N4401_1 ( .fault(fault), .net(N4401), .FEN(FEN[2617]), .op(N4401_t1) );
fim FAN_N4401_2 ( .fault(fault), .net(N4401), .FEN(FEN[2618]), .op(N4401_t2) );
fim FAN_N4405_0 ( .fault(fault), .net(N4405), .FEN(FEN[2619]), .op(N4405_t0) );
fim FAN_N4405_1 ( .fault(fault), .net(N4405), .FEN(FEN[2620]), .op(N4405_t1) );
fim FAN_N573_0 ( .fault(fault), .net(N573), .FEN(FEN[2621]), .op(N573_t0) );
fim FAN_N573_1 ( .fault(fault), .net(N573), .FEN(FEN[2622]), .op(N573_t1) );
fim FAN_N4408_0 ( .fault(fault), .net(N4408), .FEN(FEN[2623]), .op(N4408_t0) );
fim FAN_N4408_1 ( .fault(fault), .net(N4408), .FEN(FEN[2624]), .op(N4408_t1) );
fim FAN_N621_0 ( .fault(fault), .net(N621), .FEN(FEN[2625]), .op(N621_t0) );
fim FAN_N621_1 ( .fault(fault), .net(N621), .FEN(FEN[2626]), .op(N621_t1) );
fim FAN_N4411_0 ( .fault(fault), .net(N4411), .FEN(FEN[2627]), .op(N4411_t0) );
fim FAN_N4411_1 ( .fault(fault), .net(N4411), .FEN(FEN[2628]), .op(N4411_t1) );
fim FAN_N669_0 ( .fault(fault), .net(N669), .FEN(FEN[2629]), .op(N669_t0) );
fim FAN_N669_1 ( .fault(fault), .net(N669), .FEN(FEN[2630]), .op(N669_t1) );
fim FAN_N4414_0 ( .fault(fault), .net(N4414), .FEN(FEN[2631]), .op(N4414_t0) );
fim FAN_N4414_1 ( .fault(fault), .net(N4414), .FEN(FEN[2632]), .op(N4414_t1) );
fim FAN_N717_0 ( .fault(fault), .net(N717), .FEN(FEN[2633]), .op(N717_t0) );
fim FAN_N717_1 ( .fault(fault), .net(N717), .FEN(FEN[2634]), .op(N717_t1) );
fim FAN_N4417_0 ( .fault(fault), .net(N4417), .FEN(FEN[2635]), .op(N4417_t0) );
fim FAN_N4417_1 ( .fault(fault), .net(N4417), .FEN(FEN[2636]), .op(N4417_t1) );
fim FAN_N765_0 ( .fault(fault), .net(N765), .FEN(FEN[2637]), .op(N765_t0) );
fim FAN_N765_1 ( .fault(fault), .net(N765), .FEN(FEN[2638]), .op(N765_t1) );
fim FAN_N4420_0 ( .fault(fault), .net(N4420), .FEN(FEN[2639]), .op(N4420_t0) );
fim FAN_N4420_1 ( .fault(fault), .net(N4420), .FEN(FEN[2640]), .op(N4420_t1) );
fim FAN_N813_0 ( .fault(fault), .net(N813), .FEN(FEN[2641]), .op(N813_t0) );
fim FAN_N813_1 ( .fault(fault), .net(N813), .FEN(FEN[2642]), .op(N813_t1) );
fim FAN_N4423_0 ( .fault(fault), .net(N4423), .FEN(FEN[2643]), .op(N4423_t0) );
fim FAN_N4423_1 ( .fault(fault), .net(N4423), .FEN(FEN[2644]), .op(N4423_t1) );
fim FAN_N4423_2 ( .fault(fault), .net(N4423), .FEN(FEN[2645]), .op(N4423_t2) );
fim FAN_N4432_0 ( .fault(fault), .net(N4432), .FEN(FEN[2646]), .op(N4432_t0) );
fim FAN_N4432_1 ( .fault(fault), .net(N4432), .FEN(FEN[2647]), .op(N4432_t1) );
fim FAN_N4429_0 ( .fault(fault), .net(N4429), .FEN(FEN[2648]), .op(N4429_t0) );
fim FAN_N4429_1 ( .fault(fault), .net(N4429), .FEN(FEN[2649]), .op(N4429_t1) );
fim FAN_N4435_0 ( .fault(fault), .net(N4435), .FEN(FEN[2650]), .op(N4435_t0) );
fim FAN_N4435_1 ( .fault(fault), .net(N4435), .FEN(FEN[2651]), .op(N4435_t1) );
fim FAN_N4435_2 ( .fault(fault), .net(N4435), .FEN(FEN[2652]), .op(N4435_t2) );
fim FAN_N4441_0 ( .fault(fault), .net(N4441), .FEN(FEN[2653]), .op(N4441_t0) );
fim FAN_N4441_1 ( .fault(fault), .net(N4441), .FEN(FEN[2654]), .op(N4441_t1) );
fim FAN_N1056_0 ( .fault(fault), .net(N1056), .FEN(FEN[2655]), .op(N1056_t0) );
fim FAN_N1056_1 ( .fault(fault), .net(N1056), .FEN(FEN[2656]), .op(N1056_t1) );
fim FAN_N4444_0 ( .fault(fault), .net(N4444), .FEN(FEN[2657]), .op(N4444_t0) );
fim FAN_N4444_1 ( .fault(fault), .net(N4444), .FEN(FEN[2658]), .op(N4444_t1) );
fim FAN_N4444_2 ( .fault(fault), .net(N4444), .FEN(FEN[2659]), .op(N4444_t2) );
fim FAN_N4453_0 ( .fault(fault), .net(N4453), .FEN(FEN[2660]), .op(N4453_t0) );
fim FAN_N4453_1 ( .fault(fault), .net(N4453), .FEN(FEN[2661]), .op(N4453_t1) );
fim FAN_N4450_0 ( .fault(fault), .net(N4450), .FEN(FEN[2662]), .op(N4450_t0) );
fim FAN_N4450_1 ( .fault(fault), .net(N4450), .FEN(FEN[2663]), .op(N4450_t1) );
fim FAN_N4456_0 ( .fault(fault), .net(N4456), .FEN(FEN[2664]), .op(N4456_t0) );
fim FAN_N4456_1 ( .fault(fault), .net(N4456), .FEN(FEN[2665]), .op(N4456_t1) );
fim FAN_N4456_2 ( .fault(fault), .net(N4456), .FEN(FEN[2666]), .op(N4456_t2) );
fim FAN_N4462_0 ( .fault(fault), .net(N4462), .FEN(FEN[2667]), .op(N4462_t0) );
fim FAN_N4462_1 ( .fault(fault), .net(N4462), .FEN(FEN[2668]), .op(N4462_t1) );
fim FAN_N4462_2 ( .fault(fault), .net(N4462), .FEN(FEN[2669]), .op(N4462_t2) );
fim FAN_N4466_0 ( .fault(fault), .net(N4466), .FEN(FEN[2670]), .op(N4466_t0) );
fim FAN_N4466_1 ( .fault(fault), .net(N4466), .FEN(FEN[2671]), .op(N4466_t1) );
fim FAN_N4466_2 ( .fault(fault), .net(N4466), .FEN(FEN[2672]), .op(N4466_t2) );
fim FAN_N4470_0 ( .fault(fault), .net(N4470), .FEN(FEN[2673]), .op(N4470_t0) );
fim FAN_N4470_1 ( .fault(fault), .net(N4470), .FEN(FEN[2674]), .op(N4470_t1) );
fim FAN_N4470_2 ( .fault(fault), .net(N4470), .FEN(FEN[2675]), .op(N4470_t2) );
fim FAN_N4474_0 ( .fault(fault), .net(N4474), .FEN(FEN[2676]), .op(N4474_t0) );
fim FAN_N4474_1 ( .fault(fault), .net(N4474), .FEN(FEN[2677]), .op(N4474_t1) );
fim FAN_N4474_2 ( .fault(fault), .net(N4474), .FEN(FEN[2678]), .op(N4474_t2) );
fim FAN_N4478_0 ( .fault(fault), .net(N4478), .FEN(FEN[2679]), .op(N4478_t0) );
fim FAN_N4478_1 ( .fault(fault), .net(N4478), .FEN(FEN[2680]), .op(N4478_t1) );
fim FAN_N4478_2 ( .fault(fault), .net(N4478), .FEN(FEN[2681]), .op(N4478_t2) );
fim FAN_N4482_0 ( .fault(fault), .net(N4482), .FEN(FEN[2682]), .op(N4482_t0) );
fim FAN_N4482_1 ( .fault(fault), .net(N4482), .FEN(FEN[2683]), .op(N4482_t1) );
fim FAN_N4482_2 ( .fault(fault), .net(N4482), .FEN(FEN[2684]), .op(N4482_t2) );
fim FAN_N4491_0 ( .fault(fault), .net(N4491), .FEN(FEN[2685]), .op(N4491_t0) );
fim FAN_N4491_1 ( .fault(fault), .net(N4491), .FEN(FEN[2686]), .op(N4491_t1) );
fim FAN_N4488_0 ( .fault(fault), .net(N4488), .FEN(FEN[2687]), .op(N4488_t0) );
fim FAN_N4488_1 ( .fault(fault), .net(N4488), .FEN(FEN[2688]), .op(N4488_t1) );
fim FAN_N4494_0 ( .fault(fault), .net(N4494), .FEN(FEN[2689]), .op(N4494_t0) );
fim FAN_N4494_1 ( .fault(fault), .net(N4494), .FEN(FEN[2690]), .op(N4494_t1) );
fim FAN_N4494_2 ( .fault(fault), .net(N4494), .FEN(FEN[2691]), .op(N4494_t2) );
fim FAN_N4500_0 ( .fault(fault), .net(N4500), .FEN(FEN[2692]), .op(N4500_t0) );
fim FAN_N4500_1 ( .fault(fault), .net(N4500), .FEN(FEN[2693]), .op(N4500_t1) );
fim FAN_N1008_0 ( .fault(fault), .net(N1008), .FEN(FEN[2694]), .op(N1008_t0) );
fim FAN_N1008_1 ( .fault(fault), .net(N1008), .FEN(FEN[2695]), .op(N1008_t1) );
fim FAN_N4503_0 ( .fault(fault), .net(N4503), .FEN(FEN[2696]), .op(N4503_t0) );
fim FAN_N4503_1 ( .fault(fault), .net(N4503), .FEN(FEN[2697]), .op(N4503_t1) );
fim FAN_N4503_2 ( .fault(fault), .net(N4503), .FEN(FEN[2698]), .op(N4503_t2) );
fim FAN_N4512_0 ( .fault(fault), .net(N4512), .FEN(FEN[2699]), .op(N4512_t0) );
fim FAN_N4512_1 ( .fault(fault), .net(N4512), .FEN(FEN[2700]), .op(N4512_t1) );
fim FAN_N4509_0 ( .fault(fault), .net(N4509), .FEN(FEN[2701]), .op(N4509_t0) );
fim FAN_N4509_1 ( .fault(fault), .net(N4509), .FEN(FEN[2702]), .op(N4509_t1) );
fim FAN_N4515_0 ( .fault(fault), .net(N4515), .FEN(FEN[2703]), .op(N4515_t0) );
fim FAN_N4515_1 ( .fault(fault), .net(N4515), .FEN(FEN[2704]), .op(N4515_t1) );
fim FAN_N4515_2 ( .fault(fault), .net(N4515), .FEN(FEN[2705]), .op(N4515_t2) );
fim FAN_N4521_0 ( .fault(fault), .net(N4521), .FEN(FEN[2706]), .op(N4521_t0) );
fim FAN_N4521_1 ( .fault(fault), .net(N4521), .FEN(FEN[2707]), .op(N4521_t1) );
fim FAN_N1251_0 ( .fault(fault), .net(N1251), .FEN(FEN[2708]), .op(N1251_t0) );
fim FAN_N1251_1 ( .fault(fault), .net(N1251), .FEN(FEN[2709]), .op(N1251_t1) );
fim FAN_N4554_0 ( .fault(fault), .net(N4554), .FEN(FEN[2710]), .op(N4554_t0) );
fim FAN_N4554_1 ( .fault(fault), .net(N4554), .FEN(FEN[2711]), .op(N4554_t1) );
fim FAN_N4551_0 ( .fault(fault), .net(N4551), .FEN(FEN[2712]), .op(N4551_t0) );
fim FAN_N4551_1 ( .fault(fault), .net(N4551), .FEN(FEN[2713]), .op(N4551_t1) );
fim FAN_N4557_0 ( .fault(fault), .net(N4557), .FEN(FEN[2714]), .op(N4557_t0) );
fim FAN_N4557_1 ( .fault(fault), .net(N4557), .FEN(FEN[2715]), .op(N4557_t1) );
fim FAN_N4557_2 ( .fault(fault), .net(N4557), .FEN(FEN[2716]), .op(N4557_t2) );
fim FAN_N4563_0 ( .fault(fault), .net(N4563), .FEN(FEN[2717]), .op(N4563_t0) );
fim FAN_N4563_1 ( .fault(fault), .net(N4563), .FEN(FEN[2718]), .op(N4563_t1) );
fim FAN_N960_0 ( .fault(fault), .net(N960), .FEN(FEN[2719]), .op(N960_t0) );
fim FAN_N960_1 ( .fault(fault), .net(N960), .FEN(FEN[2720]), .op(N960_t1) );
fim FAN_N4566_0 ( .fault(fault), .net(N4566), .FEN(FEN[2721]), .op(N4566_t0) );
fim FAN_N4566_1 ( .fault(fault), .net(N4566), .FEN(FEN[2722]), .op(N4566_t1) );
fim FAN_N4566_2 ( .fault(fault), .net(N4566), .FEN(FEN[2723]), .op(N4566_t2) );
fim FAN_N4575_0 ( .fault(fault), .net(N4575), .FEN(FEN[2724]), .op(N4575_t0) );
fim FAN_N4575_1 ( .fault(fault), .net(N4575), .FEN(FEN[2725]), .op(N4575_t1) );
fim FAN_N4572_0 ( .fault(fault), .net(N4572), .FEN(FEN[2726]), .op(N4572_t0) );
fim FAN_N4572_1 ( .fault(fault), .net(N4572), .FEN(FEN[2727]), .op(N4572_t1) );
fim FAN_N4578_0 ( .fault(fault), .net(N4578), .FEN(FEN[2728]), .op(N4578_t0) );
fim FAN_N4578_1 ( .fault(fault), .net(N4578), .FEN(FEN[2729]), .op(N4578_t1) );
fim FAN_N4578_2 ( .fault(fault), .net(N4578), .FEN(FEN[2730]), .op(N4578_t2) );
fim FAN_N4584_0 ( .fault(fault), .net(N4584), .FEN(FEN[2731]), .op(N4584_t0) );
fim FAN_N4584_1 ( .fault(fault), .net(N4584), .FEN(FEN[2732]), .op(N4584_t1) );
fim FAN_N1203_0 ( .fault(fault), .net(N1203), .FEN(FEN[2733]), .op(N1203_t0) );
fim FAN_N1203_1 ( .fault(fault), .net(N1203), .FEN(FEN[2734]), .op(N1203_t1) );
fim FAN_N4587_0 ( .fault(fault), .net(N4587), .FEN(FEN[2735]), .op(N4587_t0) );
fim FAN_N4587_1 ( .fault(fault), .net(N4587), .FEN(FEN[2736]), .op(N4587_t1) );
fim FAN_N4587_2 ( .fault(fault), .net(N4587), .FEN(FEN[2737]), .op(N4587_t2) );
fim FAN_N4592_0 ( .fault(fault), .net(N4592), .FEN(FEN[2738]), .op(N4592_t0) );
fim FAN_N4592_1 ( .fault(fault), .net(N4592), .FEN(FEN[2739]), .op(N4592_t1) );
fim FAN_N4526_0 ( .fault(fault), .net(N4526), .FEN(FEN[2740]), .op(N4526_t0) );
fim FAN_N4526_1 ( .fault(fault), .net(N4526), .FEN(FEN[2741]), .op(N4526_t1) );
fim FAN_N4595_0 ( .fault(fault), .net(N4595), .FEN(FEN[2742]), .op(N4595_t0) );
fim FAN_N4595_1 ( .fault(fault), .net(N4595), .FEN(FEN[2743]), .op(N4595_t1) );
fim FAN_N4531_0 ( .fault(fault), .net(N4531), .FEN(FEN[2744]), .op(N4531_t0) );
fim FAN_N4531_1 ( .fault(fault), .net(N4531), .FEN(FEN[2745]), .op(N4531_t1) );
fim FAN_N4598_0 ( .fault(fault), .net(N4598), .FEN(FEN[2746]), .op(N4598_t0) );
fim FAN_N4598_1 ( .fault(fault), .net(N4598), .FEN(FEN[2747]), .op(N4598_t1) );
fim FAN_N4536_0 ( .fault(fault), .net(N4536), .FEN(FEN[2748]), .op(N4536_t0) );
fim FAN_N4536_1 ( .fault(fault), .net(N4536), .FEN(FEN[2749]), .op(N4536_t1) );
fim FAN_N4601_0 ( .fault(fault), .net(N4601), .FEN(FEN[2750]), .op(N4601_t0) );
fim FAN_N4601_1 ( .fault(fault), .net(N4601), .FEN(FEN[2751]), .op(N4601_t1) );
fim FAN_N4541_0 ( .fault(fault), .net(N4541), .FEN(FEN[2752]), .op(N4541_t0) );
fim FAN_N4541_1 ( .fault(fault), .net(N4541), .FEN(FEN[2753]), .op(N4541_t1) );
fim FAN_N4604_0 ( .fault(fault), .net(N4604), .FEN(FEN[2754]), .op(N4604_t0) );
fim FAN_N4604_1 ( .fault(fault), .net(N4604), .FEN(FEN[2755]), .op(N4604_t1) );
fim FAN_N4546_0 ( .fault(fault), .net(N4546), .FEN(FEN[2756]), .op(N4546_t0) );
fim FAN_N4546_1 ( .fault(fault), .net(N4546), .FEN(FEN[2757]), .op(N4546_t1) );
fim FAN_N4607_0 ( .fault(fault), .net(N4607), .FEN(FEN[2758]), .op(N4607_t0) );
fim FAN_N4607_1 ( .fault(fault), .net(N4607), .FEN(FEN[2759]), .op(N4607_t1) );
fim FAN_N4607_2 ( .fault(fault), .net(N4607), .FEN(FEN[2760]), .op(N4607_t2) );
fim FAN_N4613_0 ( .fault(fault), .net(N4613), .FEN(FEN[2761]), .op(N4613_t0) );
fim FAN_N4613_1 ( .fault(fault), .net(N4613), .FEN(FEN[2762]), .op(N4613_t1) );
fim FAN_N912_0 ( .fault(fault), .net(N912), .FEN(FEN[2763]), .op(N912_t0) );
fim FAN_N912_1 ( .fault(fault), .net(N912), .FEN(FEN[2764]), .op(N912_t1) );
fim FAN_N4616_0 ( .fault(fault), .net(N4616), .FEN(FEN[2765]), .op(N4616_t0) );
fim FAN_N4616_1 ( .fault(fault), .net(N4616), .FEN(FEN[2766]), .op(N4616_t1) );
fim FAN_N4616_2 ( .fault(fault), .net(N4616), .FEN(FEN[2767]), .op(N4616_t2) );
fim FAN_N4625_0 ( .fault(fault), .net(N4625), .FEN(FEN[2768]), .op(N4625_t0) );
fim FAN_N4625_1 ( .fault(fault), .net(N4625), .FEN(FEN[2769]), .op(N4625_t1) );
fim FAN_N4622_0 ( .fault(fault), .net(N4622), .FEN(FEN[2770]), .op(N4622_t0) );
fim FAN_N4622_1 ( .fault(fault), .net(N4622), .FEN(FEN[2771]), .op(N4622_t1) );
fim FAN_N4628_0 ( .fault(fault), .net(N4628), .FEN(FEN[2772]), .op(N4628_t0) );
fim FAN_N4628_1 ( .fault(fault), .net(N4628), .FEN(FEN[2773]), .op(N4628_t1) );
fim FAN_N4628_2 ( .fault(fault), .net(N4628), .FEN(FEN[2774]), .op(N4628_t2) );
fim FAN_N4634_0 ( .fault(fault), .net(N4634), .FEN(FEN[2775]), .op(N4634_t0) );
fim FAN_N4634_1 ( .fault(fault), .net(N4634), .FEN(FEN[2776]), .op(N4634_t1) );
fim FAN_N1155_0 ( .fault(fault), .net(N1155), .FEN(FEN[2777]), .op(N1155_t0) );
fim FAN_N1155_1 ( .fault(fault), .net(N1155), .FEN(FEN[2778]), .op(N1155_t1) );
fim FAN_N4637_0 ( .fault(fault), .net(N4637), .FEN(FEN[2779]), .op(N4637_t0) );
fim FAN_N4637_1 ( .fault(fault), .net(N4637), .FEN(FEN[2780]), .op(N4637_t1) );
fim FAN_N4637_2 ( .fault(fault), .net(N4637), .FEN(FEN[2781]), .op(N4637_t2) );
fim FAN_N1299_0 ( .fault(fault), .net(N1299), .FEN(FEN[2782]), .op(N1299_t0) );
fim FAN_N1299_1 ( .fault(fault), .net(N1299), .FEN(FEN[2783]), .op(N1299_t1) );
fim FAN_N4643_0 ( .fault(fault), .net(N4643), .FEN(FEN[2784]), .op(N4643_t0) );
fim FAN_N4643_1 ( .fault(fault), .net(N4643), .FEN(FEN[2785]), .op(N4643_t1) );
fim FAN_N4646_0 ( .fault(fault), .net(N4646), .FEN(FEN[2786]), .op(N4646_t0) );
fim FAN_N4646_1 ( .fault(fault), .net(N4646), .FEN(FEN[2787]), .op(N4646_t1) );
fim FAN_N4646_2 ( .fault(fault), .net(N4646), .FEN(FEN[2788]), .op(N4646_t2) );
fim FAN_N4650_0 ( .fault(fault), .net(N4650), .FEN(FEN[2789]), .op(N4650_t0) );
fim FAN_N4650_1 ( .fault(fault), .net(N4650), .FEN(FEN[2790]), .op(N4650_t1) );
fim FAN_N4650_2 ( .fault(fault), .net(N4650), .FEN(FEN[2791]), .op(N4650_t2) );
fim FAN_N4654_0 ( .fault(fault), .net(N4654), .FEN(FEN[2792]), .op(N4654_t0) );
fim FAN_N4654_1 ( .fault(fault), .net(N4654), .FEN(FEN[2793]), .op(N4654_t1) );
fim FAN_N4654_2 ( .fault(fault), .net(N4654), .FEN(FEN[2794]), .op(N4654_t2) );
fim FAN_N4658_0 ( .fault(fault), .net(N4658), .FEN(FEN[2795]), .op(N4658_t0) );
fim FAN_N4658_1 ( .fault(fault), .net(N4658), .FEN(FEN[2796]), .op(N4658_t1) );
fim FAN_N4658_2 ( .fault(fault), .net(N4658), .FEN(FEN[2797]), .op(N4658_t2) );
fim FAN_N4662_0 ( .fault(fault), .net(N4662), .FEN(FEN[2798]), .op(N4662_t0) );
fim FAN_N4662_1 ( .fault(fault), .net(N4662), .FEN(FEN[2799]), .op(N4662_t1) );
fim FAN_N4662_2 ( .fault(fault), .net(N4662), .FEN(FEN[2800]), .op(N4662_t2) );
fim FAN_N4668_0 ( .fault(fault), .net(N4668), .FEN(FEN[2801]), .op(N4668_t0) );
fim FAN_N4668_1 ( .fault(fault), .net(N4668), .FEN(FEN[2802]), .op(N4668_t1) );
fim FAN_N864_0 ( .fault(fault), .net(N864), .FEN(FEN[2803]), .op(N864_t0) );
fim FAN_N864_1 ( .fault(fault), .net(N864), .FEN(FEN[2804]), .op(N864_t1) );
fim FAN_N4671_0 ( .fault(fault), .net(N4671), .FEN(FEN[2805]), .op(N4671_t0) );
fim FAN_N4671_1 ( .fault(fault), .net(N4671), .FEN(FEN[2806]), .op(N4671_t1) );
fim FAN_N4671_2 ( .fault(fault), .net(N4671), .FEN(FEN[2807]), .op(N4671_t2) );
fim FAN_N4680_0 ( .fault(fault), .net(N4680), .FEN(FEN[2808]), .op(N4680_t0) );
fim FAN_N4680_1 ( .fault(fault), .net(N4680), .FEN(FEN[2809]), .op(N4680_t1) );
fim FAN_N4677_0 ( .fault(fault), .net(N4677), .FEN(FEN[2810]), .op(N4677_t0) );
fim FAN_N4677_1 ( .fault(fault), .net(N4677), .FEN(FEN[2811]), .op(N4677_t1) );
fim FAN_N4683_0 ( .fault(fault), .net(N4683), .FEN(FEN[2812]), .op(N4683_t0) );
fim FAN_N4683_1 ( .fault(fault), .net(N4683), .FEN(FEN[2813]), .op(N4683_t1) );
fim FAN_N4683_2 ( .fault(fault), .net(N4683), .FEN(FEN[2814]), .op(N4683_t2) );
fim FAN_N4689_0 ( .fault(fault), .net(N4689), .FEN(FEN[2815]), .op(N4689_t0) );
fim FAN_N4689_1 ( .fault(fault), .net(N4689), .FEN(FEN[2816]), .op(N4689_t1) );
fim FAN_N1107_0 ( .fault(fault), .net(N1107), .FEN(FEN[2817]), .op(N1107_t0) );
fim FAN_N1107_1 ( .fault(fault), .net(N1107), .FEN(FEN[2818]), .op(N1107_t1) );
fim FAN_N4692_0 ( .fault(fault), .net(N4692), .FEN(FEN[2819]), .op(N4692_t0) );
fim FAN_N4692_1 ( .fault(fault), .net(N4692), .FEN(FEN[2820]), .op(N4692_t1) );
fim FAN_N4692_2 ( .fault(fault), .net(N4692), .FEN(FEN[2821]), .op(N4692_t2) );
fim FAN_N4701_0 ( .fault(fault), .net(N4701), .FEN(FEN[2822]), .op(N4701_t0) );
fim FAN_N4701_1 ( .fault(fault), .net(N4701), .FEN(FEN[2823]), .op(N4701_t1) );
fim FAN_N4698_0 ( .fault(fault), .net(N4698), .FEN(FEN[2824]), .op(N4698_t0) );
fim FAN_N4698_1 ( .fault(fault), .net(N4698), .FEN(FEN[2825]), .op(N4698_t1) );
fim FAN_N4704_0 ( .fault(fault), .net(N4704), .FEN(FEN[2826]), .op(N4704_t0) );
fim FAN_N4704_1 ( .fault(fault), .net(N4704), .FEN(FEN[2827]), .op(N4704_t1) );
fim FAN_N4704_2 ( .fault(fault), .net(N4704), .FEN(FEN[2828]), .op(N4704_t2) );
fim FAN_N4718_0 ( .fault(fault), .net(N4718), .FEN(FEN[2829]), .op(N4718_t0) );
fim FAN_N4718_1 ( .fault(fault), .net(N4718), .FEN(FEN[2830]), .op(N4718_t1) );
fim FAN_N816_0 ( .fault(fault), .net(N816), .FEN(FEN[2831]), .op(N816_t0) );
fim FAN_N816_1 ( .fault(fault), .net(N816), .FEN(FEN[2832]), .op(N816_t1) );
fim FAN_N4721_0 ( .fault(fault), .net(N4721), .FEN(FEN[2833]), .op(N4721_t0) );
fim FAN_N4721_1 ( .fault(fault), .net(N4721), .FEN(FEN[2834]), .op(N4721_t1) );
fim FAN_N4721_2 ( .fault(fault), .net(N4721), .FEN(FEN[2835]), .op(N4721_t2) );
fim FAN_N4730_0 ( .fault(fault), .net(N4730), .FEN(FEN[2836]), .op(N4730_t0) );
fim FAN_N4730_1 ( .fault(fault), .net(N4730), .FEN(FEN[2837]), .op(N4730_t1) );
fim FAN_N4727_0 ( .fault(fault), .net(N4727), .FEN(FEN[2838]), .op(N4727_t0) );
fim FAN_N4727_1 ( .fault(fault), .net(N4727), .FEN(FEN[2839]), .op(N4727_t1) );
fim FAN_N4733_0 ( .fault(fault), .net(N4733), .FEN(FEN[2840]), .op(N4733_t0) );
fim FAN_N4733_1 ( .fault(fault), .net(N4733), .FEN(FEN[2841]), .op(N4733_t1) );
fim FAN_N4733_2 ( .fault(fault), .net(N4733), .FEN(FEN[2842]), .op(N4733_t2) );
fim FAN_N4739_0 ( .fault(fault), .net(N4739), .FEN(FEN[2843]), .op(N4739_t0) );
fim FAN_N4739_1 ( .fault(fault), .net(N4739), .FEN(FEN[2844]), .op(N4739_t1) );
fim FAN_N1059_0 ( .fault(fault), .net(N1059), .FEN(FEN[2845]), .op(N1059_t0) );
fim FAN_N1059_1 ( .fault(fault), .net(N1059), .FEN(FEN[2846]), .op(N1059_t1) );
fim FAN_N4742_0 ( .fault(fault), .net(N4742), .FEN(FEN[2847]), .op(N4742_t0) );
fim FAN_N4742_1 ( .fault(fault), .net(N4742), .FEN(FEN[2848]), .op(N4742_t1) );
fim FAN_N4742_2 ( .fault(fault), .net(N4742), .FEN(FEN[2849]), .op(N4742_t2) );
fim FAN_N4751_0 ( .fault(fault), .net(N4751), .FEN(FEN[2850]), .op(N4751_t0) );
fim FAN_N4751_1 ( .fault(fault), .net(N4751), .FEN(FEN[2851]), .op(N4751_t1) );
fim FAN_N4748_0 ( .fault(fault), .net(N4748), .FEN(FEN[2852]), .op(N4748_t0) );
fim FAN_N4748_1 ( .fault(fault), .net(N4748), .FEN(FEN[2853]), .op(N4748_t1) );
fim FAN_N4754_0 ( .fault(fault), .net(N4754), .FEN(FEN[2854]), .op(N4754_t0) );
fim FAN_N4754_1 ( .fault(fault), .net(N4754), .FEN(FEN[2855]), .op(N4754_t1) );
fim FAN_N4754_2 ( .fault(fault), .net(N4754), .FEN(FEN[2856]), .op(N4754_t2) );
fim FAN_N4760_0 ( .fault(fault), .net(N4760), .FEN(FEN[2857]), .op(N4760_t0) );
fim FAN_N4760_1 ( .fault(fault), .net(N4760), .FEN(FEN[2858]), .op(N4760_t1) );
fim FAN_N576_0 ( .fault(fault), .net(N576), .FEN(FEN[2859]), .op(N576_t0) );
fim FAN_N576_1 ( .fault(fault), .net(N576), .FEN(FEN[2860]), .op(N576_t1) );
fim FAN_N4763_0 ( .fault(fault), .net(N4763), .FEN(FEN[2861]), .op(N4763_t0) );
fim FAN_N4763_1 ( .fault(fault), .net(N4763), .FEN(FEN[2862]), .op(N4763_t1) );
fim FAN_N624_0 ( .fault(fault), .net(N624), .FEN(FEN[2863]), .op(N624_t0) );
fim FAN_N624_1 ( .fault(fault), .net(N624), .FEN(FEN[2864]), .op(N624_t1) );
fim FAN_N4766_0 ( .fault(fault), .net(N4766), .FEN(FEN[2865]), .op(N4766_t0) );
fim FAN_N4766_1 ( .fault(fault), .net(N4766), .FEN(FEN[2866]), .op(N4766_t1) );
fim FAN_N672_0 ( .fault(fault), .net(N672), .FEN(FEN[2867]), .op(N672_t0) );
fim FAN_N672_1 ( .fault(fault), .net(N672), .FEN(FEN[2868]), .op(N672_t1) );
fim FAN_N4769_0 ( .fault(fault), .net(N4769), .FEN(FEN[2869]), .op(N4769_t0) );
fim FAN_N4769_1 ( .fault(fault), .net(N4769), .FEN(FEN[2870]), .op(N4769_t1) );
fim FAN_N720_0 ( .fault(fault), .net(N720), .FEN(FEN[2871]), .op(N720_t0) );
fim FAN_N720_1 ( .fault(fault), .net(N720), .FEN(FEN[2872]), .op(N720_t1) );
fim FAN_N4772_0 ( .fault(fault), .net(N4772), .FEN(FEN[2873]), .op(N4772_t0) );
fim FAN_N4772_1 ( .fault(fault), .net(N4772), .FEN(FEN[2874]), .op(N4772_t1) );
fim FAN_N768_0 ( .fault(fault), .net(N768), .FEN(FEN[2875]), .op(N768_t0) );
fim FAN_N768_1 ( .fault(fault), .net(N768), .FEN(FEN[2876]), .op(N768_t1) );
fim FAN_N4775_0 ( .fault(fault), .net(N4775), .FEN(FEN[2877]), .op(N4775_t0) );
fim FAN_N4775_1 ( .fault(fault), .net(N4775), .FEN(FEN[2878]), .op(N4775_t1) );
fim FAN_N4775_2 ( .fault(fault), .net(N4775), .FEN(FEN[2879]), .op(N4775_t2) );
fim FAN_N4784_0 ( .fault(fault), .net(N4784), .FEN(FEN[2880]), .op(N4784_t0) );
fim FAN_N4784_1 ( .fault(fault), .net(N4784), .FEN(FEN[2881]), .op(N4784_t1) );
fim FAN_N4781_0 ( .fault(fault), .net(N4781), .FEN(FEN[2882]), .op(N4781_t0) );
fim FAN_N4781_1 ( .fault(fault), .net(N4781), .FEN(FEN[2883]), .op(N4781_t1) );
fim FAN_N4787_0 ( .fault(fault), .net(N4787), .FEN(FEN[2884]), .op(N4787_t0) );
fim FAN_N4787_1 ( .fault(fault), .net(N4787), .FEN(FEN[2885]), .op(N4787_t1) );
fim FAN_N4787_2 ( .fault(fault), .net(N4787), .FEN(FEN[2886]), .op(N4787_t2) );
fim FAN_N4793_0 ( .fault(fault), .net(N4793), .FEN(FEN[2887]), .op(N4793_t0) );
fim FAN_N4793_1 ( .fault(fault), .net(N4793), .FEN(FEN[2888]), .op(N4793_t1) );
fim FAN_N1011_0 ( .fault(fault), .net(N1011), .FEN(FEN[2889]), .op(N1011_t0) );
fim FAN_N1011_1 ( .fault(fault), .net(N1011), .FEN(FEN[2890]), .op(N1011_t1) );
fim FAN_N4796_0 ( .fault(fault), .net(N4796), .FEN(FEN[2891]), .op(N4796_t0) );
fim FAN_N4796_1 ( .fault(fault), .net(N4796), .FEN(FEN[2892]), .op(N4796_t1) );
fim FAN_N4796_2 ( .fault(fault), .net(N4796), .FEN(FEN[2893]), .op(N4796_t2) );
fim FAN_N4805_0 ( .fault(fault), .net(N4805), .FEN(FEN[2894]), .op(N4805_t0) );
fim FAN_N4805_1 ( .fault(fault), .net(N4805), .FEN(FEN[2895]), .op(N4805_t1) );
fim FAN_N4802_0 ( .fault(fault), .net(N4802), .FEN(FEN[2896]), .op(N4802_t0) );
fim FAN_N4802_1 ( .fault(fault), .net(N4802), .FEN(FEN[2897]), .op(N4802_t1) );
fim FAN_N4808_0 ( .fault(fault), .net(N4808), .FEN(FEN[2898]), .op(N4808_t0) );
fim FAN_N4808_1 ( .fault(fault), .net(N4808), .FEN(FEN[2899]), .op(N4808_t1) );
fim FAN_N4808_2 ( .fault(fault), .net(N4808), .FEN(FEN[2900]), .op(N4808_t2) );
fim FAN_N4814_0 ( .fault(fault), .net(N4814), .FEN(FEN[2901]), .op(N4814_t0) );
fim FAN_N4814_1 ( .fault(fault), .net(N4814), .FEN(FEN[2902]), .op(N4814_t1) );
fim FAN_N1254_0 ( .fault(fault), .net(N1254), .FEN(FEN[2903]), .op(N1254_t0) );
fim FAN_N1254_1 ( .fault(fault), .net(N1254), .FEN(FEN[2904]), .op(N1254_t1) );
fim FAN_N4817_0 ( .fault(fault), .net(N4817), .FEN(FEN[2905]), .op(N4817_t0) );
fim FAN_N4817_1 ( .fault(fault), .net(N4817), .FEN(FEN[2906]), .op(N4817_t1) );
fim FAN_N4817_2 ( .fault(fault), .net(N4817), .FEN(FEN[2907]), .op(N4817_t2) );
fim FAN_N4821_0 ( .fault(fault), .net(N4821), .FEN(FEN[2908]), .op(N4821_t0) );
fim FAN_N4821_1 ( .fault(fault), .net(N4821), .FEN(FEN[2909]), .op(N4821_t1) );
fim FAN_N4821_2 ( .fault(fault), .net(N4821), .FEN(FEN[2910]), .op(N4821_t2) );
fim FAN_N4825_0 ( .fault(fault), .net(N4825), .FEN(FEN[2911]), .op(N4825_t0) );
fim FAN_N4825_1 ( .fault(fault), .net(N4825), .FEN(FEN[2912]), .op(N4825_t1) );
fim FAN_N4825_2 ( .fault(fault), .net(N4825), .FEN(FEN[2913]), .op(N4825_t2) );
fim FAN_N4829_0 ( .fault(fault), .net(N4829), .FEN(FEN[2914]), .op(N4829_t0) );
fim FAN_N4829_1 ( .fault(fault), .net(N4829), .FEN(FEN[2915]), .op(N4829_t1) );
fim FAN_N4829_2 ( .fault(fault), .net(N4829), .FEN(FEN[2916]), .op(N4829_t2) );
fim FAN_N4833_0 ( .fault(fault), .net(N4833), .FEN(FEN[2917]), .op(N4833_t0) );
fim FAN_N4833_1 ( .fault(fault), .net(N4833), .FEN(FEN[2918]), .op(N4833_t1) );
fim FAN_N4833_2 ( .fault(fault), .net(N4833), .FEN(FEN[2919]), .op(N4833_t2) );
fim FAN_N4842_0 ( .fault(fault), .net(N4842), .FEN(FEN[2920]), .op(N4842_t0) );
fim FAN_N4842_1 ( .fault(fault), .net(N4842), .FEN(FEN[2921]), .op(N4842_t1) );
fim FAN_N4839_0 ( .fault(fault), .net(N4839), .FEN(FEN[2922]), .op(N4839_t0) );
fim FAN_N4839_1 ( .fault(fault), .net(N4839), .FEN(FEN[2923]), .op(N4839_t1) );
fim FAN_N4845_0 ( .fault(fault), .net(N4845), .FEN(FEN[2924]), .op(N4845_t0) );
fim FAN_N4845_1 ( .fault(fault), .net(N4845), .FEN(FEN[2925]), .op(N4845_t1) );
fim FAN_N4845_2 ( .fault(fault), .net(N4845), .FEN(FEN[2926]), .op(N4845_t2) );
fim FAN_N4851_0 ( .fault(fault), .net(N4851), .FEN(FEN[2927]), .op(N4851_t0) );
fim FAN_N4851_1 ( .fault(fault), .net(N4851), .FEN(FEN[2928]), .op(N4851_t1) );
fim FAN_N963_0 ( .fault(fault), .net(N963), .FEN(FEN[2929]), .op(N963_t0) );
fim FAN_N963_1 ( .fault(fault), .net(N963), .FEN(FEN[2930]), .op(N963_t1) );
fim FAN_N4854_0 ( .fault(fault), .net(N4854), .FEN(FEN[2931]), .op(N4854_t0) );
fim FAN_N4854_1 ( .fault(fault), .net(N4854), .FEN(FEN[2932]), .op(N4854_t1) );
fim FAN_N4854_2 ( .fault(fault), .net(N4854), .FEN(FEN[2933]), .op(N4854_t2) );
fim FAN_N4863_0 ( .fault(fault), .net(N4863), .FEN(FEN[2934]), .op(N4863_t0) );
fim FAN_N4863_1 ( .fault(fault), .net(N4863), .FEN(FEN[2935]), .op(N4863_t1) );
fim FAN_N4860_0 ( .fault(fault), .net(N4860), .FEN(FEN[2936]), .op(N4860_t0) );
fim FAN_N4860_1 ( .fault(fault), .net(N4860), .FEN(FEN[2937]), .op(N4860_t1) );
fim FAN_N4866_0 ( .fault(fault), .net(N4866), .FEN(FEN[2938]), .op(N4866_t0) );
fim FAN_N4866_1 ( .fault(fault), .net(N4866), .FEN(FEN[2939]), .op(N4866_t1) );
fim FAN_N4866_2 ( .fault(fault), .net(N4866), .FEN(FEN[2940]), .op(N4866_t2) );
fim FAN_N4872_0 ( .fault(fault), .net(N4872), .FEN(FEN[2941]), .op(N4872_t0) );
fim FAN_N4872_1 ( .fault(fault), .net(N4872), .FEN(FEN[2942]), .op(N4872_t1) );
fim FAN_N1206_0 ( .fault(fault), .net(N1206), .FEN(FEN[2943]), .op(N1206_t0) );
fim FAN_N1206_1 ( .fault(fault), .net(N1206), .FEN(FEN[2944]), .op(N1206_t1) );
fim FAN_N4875_0 ( .fault(fault), .net(N4875), .FEN(FEN[2945]), .op(N4875_t0) );
fim FAN_N4875_1 ( .fault(fault), .net(N4875), .FEN(FEN[2946]), .op(N4875_t1) );
fim FAN_N4875_2 ( .fault(fault), .net(N4875), .FEN(FEN[2947]), .op(N4875_t2) );
fim FAN_N4904_0 ( .fault(fault), .net(N4904), .FEN(FEN[2948]), .op(N4904_t0) );
fim FAN_N4904_1 ( .fault(fault), .net(N4904), .FEN(FEN[2949]), .op(N4904_t1) );
fim FAN_N4901_0 ( .fault(fault), .net(N4901), .FEN(FEN[2950]), .op(N4901_t0) );
fim FAN_N4901_1 ( .fault(fault), .net(N4901), .FEN(FEN[2951]), .op(N4901_t1) );
fim FAN_N4907_0 ( .fault(fault), .net(N4907), .FEN(FEN[2952]), .op(N4907_t0) );
fim FAN_N4907_1 ( .fault(fault), .net(N4907), .FEN(FEN[2953]), .op(N4907_t1) );
fim FAN_N4907_2 ( .fault(fault), .net(N4907), .FEN(FEN[2954]), .op(N4907_t2) );
fim FAN_N4913_0 ( .fault(fault), .net(N4913), .FEN(FEN[2955]), .op(N4913_t0) );
fim FAN_N4913_1 ( .fault(fault), .net(N4913), .FEN(FEN[2956]), .op(N4913_t1) );
fim FAN_N915_0 ( .fault(fault), .net(N915), .FEN(FEN[2957]), .op(N915_t0) );
fim FAN_N915_1 ( .fault(fault), .net(N915), .FEN(FEN[2958]), .op(N915_t1) );
fim FAN_N4916_0 ( .fault(fault), .net(N4916), .FEN(FEN[2959]), .op(N4916_t0) );
fim FAN_N4916_1 ( .fault(fault), .net(N4916), .FEN(FEN[2960]), .op(N4916_t1) );
fim FAN_N4916_2 ( .fault(fault), .net(N4916), .FEN(FEN[2961]), .op(N4916_t2) );
fim FAN_N4925_0 ( .fault(fault), .net(N4925), .FEN(FEN[2962]), .op(N4925_t0) );
fim FAN_N4925_1 ( .fault(fault), .net(N4925), .FEN(FEN[2963]), .op(N4925_t1) );
fim FAN_N4922_0 ( .fault(fault), .net(N4922), .FEN(FEN[2964]), .op(N4922_t0) );
fim FAN_N4922_1 ( .fault(fault), .net(N4922), .FEN(FEN[2965]), .op(N4922_t1) );
fim FAN_N4928_0 ( .fault(fault), .net(N4928), .FEN(FEN[2966]), .op(N4928_t0) );
fim FAN_N4928_1 ( .fault(fault), .net(N4928), .FEN(FEN[2967]), .op(N4928_t1) );
fim FAN_N4928_2 ( .fault(fault), .net(N4928), .FEN(FEN[2968]), .op(N4928_t2) );
fim FAN_N4934_0 ( .fault(fault), .net(N4934), .FEN(FEN[2969]), .op(N4934_t0) );
fim FAN_N4934_1 ( .fault(fault), .net(N4934), .FEN(FEN[2970]), .op(N4934_t1) );
fim FAN_N1158_0 ( .fault(fault), .net(N1158), .FEN(FEN[2971]), .op(N1158_t0) );
fim FAN_N1158_1 ( .fault(fault), .net(N1158), .FEN(FEN[2972]), .op(N1158_t1) );
fim FAN_N4937_0 ( .fault(fault), .net(N4937), .FEN(FEN[2973]), .op(N4937_t0) );
fim FAN_N4937_1 ( .fault(fault), .net(N4937), .FEN(FEN[2974]), .op(N4937_t1) );
fim FAN_N4937_2 ( .fault(fault), .net(N4937), .FEN(FEN[2975]), .op(N4937_t2) );
fim FAN_N1302_0 ( .fault(fault), .net(N1302), .FEN(FEN[2976]), .op(N1302_t0) );
fim FAN_N1302_1 ( .fault(fault), .net(N1302), .FEN(FEN[2977]), .op(N1302_t1) );
fim FAN_N4943_0 ( .fault(fault), .net(N4943), .FEN(FEN[2978]), .op(N4943_t0) );
fim FAN_N4943_1 ( .fault(fault), .net(N4943), .FEN(FEN[2979]), .op(N4943_t1) );
fim FAN_N4947_0 ( .fault(fault), .net(N4947), .FEN(FEN[2980]), .op(N4947_t0) );
fim FAN_N4947_1 ( .fault(fault), .net(N4947), .FEN(FEN[2981]), .op(N4947_t1) );
fim FAN_N4881_0 ( .fault(fault), .net(N4881), .FEN(FEN[2982]), .op(N4881_t0) );
fim FAN_N4881_1 ( .fault(fault), .net(N4881), .FEN(FEN[2983]), .op(N4881_t1) );
fim FAN_N4950_0 ( .fault(fault), .net(N4950), .FEN(FEN[2984]), .op(N4950_t0) );
fim FAN_N4950_1 ( .fault(fault), .net(N4950), .FEN(FEN[2985]), .op(N4950_t1) );
fim FAN_N4886_0 ( .fault(fault), .net(N4886), .FEN(FEN[2986]), .op(N4886_t0) );
fim FAN_N4886_1 ( .fault(fault), .net(N4886), .FEN(FEN[2987]), .op(N4886_t1) );
fim FAN_N4953_0 ( .fault(fault), .net(N4953), .FEN(FEN[2988]), .op(N4953_t0) );
fim FAN_N4953_1 ( .fault(fault), .net(N4953), .FEN(FEN[2989]), .op(N4953_t1) );
fim FAN_N4891_0 ( .fault(fault), .net(N4891), .FEN(FEN[2990]), .op(N4891_t0) );
fim FAN_N4891_1 ( .fault(fault), .net(N4891), .FEN(FEN[2991]), .op(N4891_t1) );
fim FAN_N4956_0 ( .fault(fault), .net(N4956), .FEN(FEN[2992]), .op(N4956_t0) );
fim FAN_N4956_1 ( .fault(fault), .net(N4956), .FEN(FEN[2993]), .op(N4956_t1) );
fim FAN_N4896_0 ( .fault(fault), .net(N4896), .FEN(FEN[2994]), .op(N4896_t0) );
fim FAN_N4896_1 ( .fault(fault), .net(N4896), .FEN(FEN[2995]), .op(N4896_t1) );
fim FAN_N4959_0 ( .fault(fault), .net(N4959), .FEN(FEN[2996]), .op(N4959_t0) );
fim FAN_N4959_1 ( .fault(fault), .net(N4959), .FEN(FEN[2997]), .op(N4959_t1) );
fim FAN_N4959_2 ( .fault(fault), .net(N4959), .FEN(FEN[2998]), .op(N4959_t2) );
fim FAN_N4965_0 ( .fault(fault), .net(N4965), .FEN(FEN[2999]), .op(N4965_t0) );
fim FAN_N4965_1 ( .fault(fault), .net(N4965), .FEN(FEN[3000]), .op(N4965_t1) );
fim FAN_N867_0 ( .fault(fault), .net(N867), .FEN(FEN[3001]), .op(N867_t0) );
fim FAN_N867_1 ( .fault(fault), .net(N867), .FEN(FEN[3002]), .op(N867_t1) );
fim FAN_N4968_0 ( .fault(fault), .net(N4968), .FEN(FEN[3003]), .op(N4968_t0) );
fim FAN_N4968_1 ( .fault(fault), .net(N4968), .FEN(FEN[3004]), .op(N4968_t1) );
fim FAN_N4968_2 ( .fault(fault), .net(N4968), .FEN(FEN[3005]), .op(N4968_t2) );
fim FAN_N4977_0 ( .fault(fault), .net(N4977), .FEN(FEN[3006]), .op(N4977_t0) );
fim FAN_N4977_1 ( .fault(fault), .net(N4977), .FEN(FEN[3007]), .op(N4977_t1) );
fim FAN_N4974_0 ( .fault(fault), .net(N4974), .FEN(FEN[3008]), .op(N4974_t0) );
fim FAN_N4974_1 ( .fault(fault), .net(N4974), .FEN(FEN[3009]), .op(N4974_t1) );
fim FAN_N4980_0 ( .fault(fault), .net(N4980), .FEN(FEN[3010]), .op(N4980_t0) );
fim FAN_N4980_1 ( .fault(fault), .net(N4980), .FEN(FEN[3011]), .op(N4980_t1) );
fim FAN_N4980_2 ( .fault(fault), .net(N4980), .FEN(FEN[3012]), .op(N4980_t2) );
fim FAN_N4986_0 ( .fault(fault), .net(N4986), .FEN(FEN[3013]), .op(N4986_t0) );
fim FAN_N4986_1 ( .fault(fault), .net(N4986), .FEN(FEN[3014]), .op(N4986_t1) );
fim FAN_N1110_0 ( .fault(fault), .net(N1110), .FEN(FEN[3015]), .op(N1110_t0) );
fim FAN_N1110_1 ( .fault(fault), .net(N1110), .FEN(FEN[3016]), .op(N1110_t1) );
fim FAN_N4989_0 ( .fault(fault), .net(N4989), .FEN(FEN[3017]), .op(N4989_t0) );
fim FAN_N4989_1 ( .fault(fault), .net(N4989), .FEN(FEN[3018]), .op(N4989_t1) );
fim FAN_N4989_2 ( .fault(fault), .net(N4989), .FEN(FEN[3019]), .op(N4989_t2) );
fim FAN_N4998_0 ( .fault(fault), .net(N4998), .FEN(FEN[3020]), .op(N4998_t0) );
fim FAN_N4998_1 ( .fault(fault), .net(N4998), .FEN(FEN[3021]), .op(N4998_t1) );
fim FAN_N4995_0 ( .fault(fault), .net(N4995), .FEN(FEN[3022]), .op(N4995_t0) );
fim FAN_N4995_1 ( .fault(fault), .net(N4995), .FEN(FEN[3023]), .op(N4995_t1) );
fim FAN_N5001_0 ( .fault(fault), .net(N5001), .FEN(FEN[3024]), .op(N5001_t0) );
fim FAN_N5001_1 ( .fault(fault), .net(N5001), .FEN(FEN[3025]), .op(N5001_t1) );
fim FAN_N5001_2 ( .fault(fault), .net(N5001), .FEN(FEN[3026]), .op(N5001_t2) );
fim FAN_N5005_0 ( .fault(fault), .net(N5005), .FEN(FEN[3027]), .op(N5005_t0) );
fim FAN_N5005_1 ( .fault(fault), .net(N5005), .FEN(FEN[3028]), .op(N5005_t1) );
fim FAN_N5005_2 ( .fault(fault), .net(N5005), .FEN(FEN[3029]), .op(N5005_t2) );
fim FAN_N5009_0 ( .fault(fault), .net(N5009), .FEN(FEN[3030]), .op(N5009_t0) );
fim FAN_N5009_1 ( .fault(fault), .net(N5009), .FEN(FEN[3031]), .op(N5009_t1) );
fim FAN_N5009_2 ( .fault(fault), .net(N5009), .FEN(FEN[3032]), .op(N5009_t2) );
fim FAN_N5013_0 ( .fault(fault), .net(N5013), .FEN(FEN[3033]), .op(N5013_t0) );
fim FAN_N5013_1 ( .fault(fault), .net(N5013), .FEN(FEN[3034]), .op(N5013_t1) );
fim FAN_N5013_2 ( .fault(fault), .net(N5013), .FEN(FEN[3035]), .op(N5013_t2) );
fim FAN_N5017_0 ( .fault(fault), .net(N5017), .FEN(FEN[3036]), .op(N5017_t0) );
fim FAN_N5017_1 ( .fault(fault), .net(N5017), .FEN(FEN[3037]), .op(N5017_t1) );
fim FAN_N5017_2 ( .fault(fault), .net(N5017), .FEN(FEN[3038]), .op(N5017_t2) );
fim FAN_N5023_0 ( .fault(fault), .net(N5023), .FEN(FEN[3039]), .op(N5023_t0) );
fim FAN_N5023_1 ( .fault(fault), .net(N5023), .FEN(FEN[3040]), .op(N5023_t1) );
fim FAN_N819_0 ( .fault(fault), .net(N819), .FEN(FEN[3041]), .op(N819_t0) );
fim FAN_N819_1 ( .fault(fault), .net(N819), .FEN(FEN[3042]), .op(N819_t1) );
fim FAN_N5026_0 ( .fault(fault), .net(N5026), .FEN(FEN[3043]), .op(N5026_t0) );
fim FAN_N5026_1 ( .fault(fault), .net(N5026), .FEN(FEN[3044]), .op(N5026_t1) );
fim FAN_N5026_2 ( .fault(fault), .net(N5026), .FEN(FEN[3045]), .op(N5026_t2) );
fim FAN_N5035_0 ( .fault(fault), .net(N5035), .FEN(FEN[3046]), .op(N5035_t0) );
fim FAN_N5035_1 ( .fault(fault), .net(N5035), .FEN(FEN[3047]), .op(N5035_t1) );
fim FAN_N5032_0 ( .fault(fault), .net(N5032), .FEN(FEN[3048]), .op(N5032_t0) );
fim FAN_N5032_1 ( .fault(fault), .net(N5032), .FEN(FEN[3049]), .op(N5032_t1) );
fim FAN_N5038_0 ( .fault(fault), .net(N5038), .FEN(FEN[3050]), .op(N5038_t0) );
fim FAN_N5038_1 ( .fault(fault), .net(N5038), .FEN(FEN[3051]), .op(N5038_t1) );
fim FAN_N5038_2 ( .fault(fault), .net(N5038), .FEN(FEN[3052]), .op(N5038_t2) );
fim FAN_N5044_0 ( .fault(fault), .net(N5044), .FEN(FEN[3053]), .op(N5044_t0) );
fim FAN_N5044_1 ( .fault(fault), .net(N5044), .FEN(FEN[3054]), .op(N5044_t1) );
fim FAN_N1062_0 ( .fault(fault), .net(N1062), .FEN(FEN[3055]), .op(N1062_t0) );
fim FAN_N1062_1 ( .fault(fault), .net(N1062), .FEN(FEN[3056]), .op(N1062_t1) );
fim FAN_N5047_0 ( .fault(fault), .net(N5047), .FEN(FEN[3057]), .op(N5047_t0) );
fim FAN_N5047_1 ( .fault(fault), .net(N5047), .FEN(FEN[3058]), .op(N5047_t1) );
fim FAN_N5047_2 ( .fault(fault), .net(N5047), .FEN(FEN[3059]), .op(N5047_t2) );
fim FAN_N5056_0 ( .fault(fault), .net(N5056), .FEN(FEN[3060]), .op(N5056_t0) );
fim FAN_N5056_1 ( .fault(fault), .net(N5056), .FEN(FEN[3061]), .op(N5056_t1) );
fim FAN_N5053_0 ( .fault(fault), .net(N5053), .FEN(FEN[3062]), .op(N5053_t0) );
fim FAN_N5053_1 ( .fault(fault), .net(N5053), .FEN(FEN[3063]), .op(N5053_t1) );
fim FAN_N5059_0 ( .fault(fault), .net(N5059), .FEN(FEN[3064]), .op(N5059_t0) );
fim FAN_N5059_1 ( .fault(fault), .net(N5059), .FEN(FEN[3065]), .op(N5059_t1) );
fim FAN_N5059_2 ( .fault(fault), .net(N5059), .FEN(FEN[3066]), .op(N5059_t2) );
fim FAN_N5073_0 ( .fault(fault), .net(N5073), .FEN(FEN[3067]), .op(N5073_t0) );
fim FAN_N5073_1 ( .fault(fault), .net(N5073), .FEN(FEN[3068]), .op(N5073_t1) );
fim FAN_N771_0 ( .fault(fault), .net(N771), .FEN(FEN[3069]), .op(N771_t0) );
fim FAN_N771_1 ( .fault(fault), .net(N771), .FEN(FEN[3070]), .op(N771_t1) );
fim FAN_N5076_0 ( .fault(fault), .net(N5076), .FEN(FEN[3071]), .op(N5076_t0) );
fim FAN_N5076_1 ( .fault(fault), .net(N5076), .FEN(FEN[3072]), .op(N5076_t1) );
fim FAN_N5076_2 ( .fault(fault), .net(N5076), .FEN(FEN[3073]), .op(N5076_t2) );
fim FAN_N5085_0 ( .fault(fault), .net(N5085), .FEN(FEN[3074]), .op(N5085_t0) );
fim FAN_N5085_1 ( .fault(fault), .net(N5085), .FEN(FEN[3075]), .op(N5085_t1) );
fim FAN_N5082_0 ( .fault(fault), .net(N5082), .FEN(FEN[3076]), .op(N5082_t0) );
fim FAN_N5082_1 ( .fault(fault), .net(N5082), .FEN(FEN[3077]), .op(N5082_t1) );
fim FAN_N5088_0 ( .fault(fault), .net(N5088), .FEN(FEN[3078]), .op(N5088_t0) );
fim FAN_N5088_1 ( .fault(fault), .net(N5088), .FEN(FEN[3079]), .op(N5088_t1) );
fim FAN_N5088_2 ( .fault(fault), .net(N5088), .FEN(FEN[3080]), .op(N5088_t2) );
fim FAN_N5094_0 ( .fault(fault), .net(N5094), .FEN(FEN[3081]), .op(N5094_t0) );
fim FAN_N5094_1 ( .fault(fault), .net(N5094), .FEN(FEN[3082]), .op(N5094_t1) );
fim FAN_N1014_0 ( .fault(fault), .net(N1014), .FEN(FEN[3083]), .op(N1014_t0) );
fim FAN_N1014_1 ( .fault(fault), .net(N1014), .FEN(FEN[3084]), .op(N1014_t1) );
fim FAN_N5097_0 ( .fault(fault), .net(N5097), .FEN(FEN[3085]), .op(N5097_t0) );
fim FAN_N5097_1 ( .fault(fault), .net(N5097), .FEN(FEN[3086]), .op(N5097_t1) );
fim FAN_N5097_2 ( .fault(fault), .net(N5097), .FEN(FEN[3087]), .op(N5097_t2) );
fim FAN_N5106_0 ( .fault(fault), .net(N5106), .FEN(FEN[3088]), .op(N5106_t0) );
fim FAN_N5106_1 ( .fault(fault), .net(N5106), .FEN(FEN[3089]), .op(N5106_t1) );
fim FAN_N5103_0 ( .fault(fault), .net(N5103), .FEN(FEN[3090]), .op(N5103_t0) );
fim FAN_N5103_1 ( .fault(fault), .net(N5103), .FEN(FEN[3091]), .op(N5103_t1) );
fim FAN_N5109_0 ( .fault(fault), .net(N5109), .FEN(FEN[3092]), .op(N5109_t0) );
fim FAN_N5109_1 ( .fault(fault), .net(N5109), .FEN(FEN[3093]), .op(N5109_t1) );
fim FAN_N5109_2 ( .fault(fault), .net(N5109), .FEN(FEN[3094]), .op(N5109_t2) );
fim FAN_N5115_0 ( .fault(fault), .net(N5115), .FEN(FEN[3095]), .op(N5115_t0) );
fim FAN_N5115_1 ( .fault(fault), .net(N5115), .FEN(FEN[3096]), .op(N5115_t1) );
fim FAN_N1257_0 ( .fault(fault), .net(N1257), .FEN(FEN[3097]), .op(N1257_t0) );
fim FAN_N1257_1 ( .fault(fault), .net(N1257), .FEN(FEN[3098]), .op(N1257_t1) );
fim FAN_N5118_0 ( .fault(fault), .net(N5118), .FEN(FEN[3099]), .op(N5118_t0) );
fim FAN_N5118_1 ( .fault(fault), .net(N5118), .FEN(FEN[3100]), .op(N5118_t1) );
fim FAN_N579_0 ( .fault(fault), .net(N579), .FEN(FEN[3101]), .op(N579_t0) );
fim FAN_N579_1 ( .fault(fault), .net(N579), .FEN(FEN[3102]), .op(N579_t1) );
fim FAN_N5121_0 ( .fault(fault), .net(N5121), .FEN(FEN[3103]), .op(N5121_t0) );
fim FAN_N5121_1 ( .fault(fault), .net(N5121), .FEN(FEN[3104]), .op(N5121_t1) );
fim FAN_N627_0 ( .fault(fault), .net(N627), .FEN(FEN[3105]), .op(N627_t0) );
fim FAN_N627_1 ( .fault(fault), .net(N627), .FEN(FEN[3106]), .op(N627_t1) );
fim FAN_N5124_0 ( .fault(fault), .net(N5124), .FEN(FEN[3107]), .op(N5124_t0) );
fim FAN_N5124_1 ( .fault(fault), .net(N5124), .FEN(FEN[3108]), .op(N5124_t1) );
fim FAN_N675_0 ( .fault(fault), .net(N675), .FEN(FEN[3109]), .op(N675_t0) );
fim FAN_N675_1 ( .fault(fault), .net(N675), .FEN(FEN[3110]), .op(N675_t1) );
fim FAN_N5127_0 ( .fault(fault), .net(N5127), .FEN(FEN[3111]), .op(N5127_t0) );
fim FAN_N5127_1 ( .fault(fault), .net(N5127), .FEN(FEN[3112]), .op(N5127_t1) );
fim FAN_N723_0 ( .fault(fault), .net(N723), .FEN(FEN[3113]), .op(N723_t0) );
fim FAN_N723_1 ( .fault(fault), .net(N723), .FEN(FEN[3114]), .op(N723_t1) );
fim FAN_N5130_0 ( .fault(fault), .net(N5130), .FEN(FEN[3115]), .op(N5130_t0) );
fim FAN_N5130_1 ( .fault(fault), .net(N5130), .FEN(FEN[3116]), .op(N5130_t1) );
fim FAN_N5130_2 ( .fault(fault), .net(N5130), .FEN(FEN[3117]), .op(N5130_t2) );
fim FAN_N5139_0 ( .fault(fault), .net(N5139), .FEN(FEN[3118]), .op(N5139_t0) );
fim FAN_N5139_1 ( .fault(fault), .net(N5139), .FEN(FEN[3119]), .op(N5139_t1) );
fim FAN_N5136_0 ( .fault(fault), .net(N5136), .FEN(FEN[3120]), .op(N5136_t0) );
fim FAN_N5136_1 ( .fault(fault), .net(N5136), .FEN(FEN[3121]), .op(N5136_t1) );
fim FAN_N5142_0 ( .fault(fault), .net(N5142), .FEN(FEN[3122]), .op(N5142_t0) );
fim FAN_N5142_1 ( .fault(fault), .net(N5142), .FEN(FEN[3123]), .op(N5142_t1) );
fim FAN_N5142_2 ( .fault(fault), .net(N5142), .FEN(FEN[3124]), .op(N5142_t2) );
fim FAN_N5148_0 ( .fault(fault), .net(N5148), .FEN(FEN[3125]), .op(N5148_t0) );
fim FAN_N5148_1 ( .fault(fault), .net(N5148), .FEN(FEN[3126]), .op(N5148_t1) );
fim FAN_N966_0 ( .fault(fault), .net(N966), .FEN(FEN[3127]), .op(N966_t0) );
fim FAN_N966_1 ( .fault(fault), .net(N966), .FEN(FEN[3128]), .op(N966_t1) );
fim FAN_N5151_0 ( .fault(fault), .net(N5151), .FEN(FEN[3129]), .op(N5151_t0) );
fim FAN_N5151_1 ( .fault(fault), .net(N5151), .FEN(FEN[3130]), .op(N5151_t1) );
fim FAN_N5151_2 ( .fault(fault), .net(N5151), .FEN(FEN[3131]), .op(N5151_t2) );
fim FAN_N5160_0 ( .fault(fault), .net(N5160), .FEN(FEN[3132]), .op(N5160_t0) );
fim FAN_N5160_1 ( .fault(fault), .net(N5160), .FEN(FEN[3133]), .op(N5160_t1) );
fim FAN_N5157_0 ( .fault(fault), .net(N5157), .FEN(FEN[3134]), .op(N5157_t0) );
fim FAN_N5157_1 ( .fault(fault), .net(N5157), .FEN(FEN[3135]), .op(N5157_t1) );
fim FAN_N5163_0 ( .fault(fault), .net(N5163), .FEN(FEN[3136]), .op(N5163_t0) );
fim FAN_N5163_1 ( .fault(fault), .net(N5163), .FEN(FEN[3137]), .op(N5163_t1) );
fim FAN_N5163_2 ( .fault(fault), .net(N5163), .FEN(FEN[3138]), .op(N5163_t2) );
fim FAN_N5169_0 ( .fault(fault), .net(N5169), .FEN(FEN[3139]), .op(N5169_t0) );
fim FAN_N5169_1 ( .fault(fault), .net(N5169), .FEN(FEN[3140]), .op(N5169_t1) );
fim FAN_N1209_0 ( .fault(fault), .net(N1209), .FEN(FEN[3141]), .op(N1209_t0) );
fim FAN_N1209_1 ( .fault(fault), .net(N1209), .FEN(FEN[3142]), .op(N1209_t1) );
fim FAN_N5172_0 ( .fault(fault), .net(N5172), .FEN(FEN[3143]), .op(N5172_t0) );
fim FAN_N5172_1 ( .fault(fault), .net(N5172), .FEN(FEN[3144]), .op(N5172_t1) );
fim FAN_N5172_2 ( .fault(fault), .net(N5172), .FEN(FEN[3145]), .op(N5172_t2) );
fim FAN_N5176_0 ( .fault(fault), .net(N5176), .FEN(FEN[3146]), .op(N5176_t0) );
fim FAN_N5176_1 ( .fault(fault), .net(N5176), .FEN(FEN[3147]), .op(N5176_t1) );
fim FAN_N5176_2 ( .fault(fault), .net(N5176), .FEN(FEN[3148]), .op(N5176_t2) );
fim FAN_N5180_0 ( .fault(fault), .net(N5180), .FEN(FEN[3149]), .op(N5180_t0) );
fim FAN_N5180_1 ( .fault(fault), .net(N5180), .FEN(FEN[3150]), .op(N5180_t1) );
fim FAN_N5180_2 ( .fault(fault), .net(N5180), .FEN(FEN[3151]), .op(N5180_t2) );
fim FAN_N5184_0 ( .fault(fault), .net(N5184), .FEN(FEN[3152]), .op(N5184_t0) );
fim FAN_N5184_1 ( .fault(fault), .net(N5184), .FEN(FEN[3153]), .op(N5184_t1) );
fim FAN_N5184_2 ( .fault(fault), .net(N5184), .FEN(FEN[3154]), .op(N5184_t2) );
fim FAN_N5188_0 ( .fault(fault), .net(N5188), .FEN(FEN[3155]), .op(N5188_t0) );
fim FAN_N5188_1 ( .fault(fault), .net(N5188), .FEN(FEN[3156]), .op(N5188_t1) );
fim FAN_N5188_2 ( .fault(fault), .net(N5188), .FEN(FEN[3157]), .op(N5188_t2) );
fim FAN_N5197_0 ( .fault(fault), .net(N5197), .FEN(FEN[3158]), .op(N5197_t0) );
fim FAN_N5197_1 ( .fault(fault), .net(N5197), .FEN(FEN[3159]), .op(N5197_t1) );
fim FAN_N5194_0 ( .fault(fault), .net(N5194), .FEN(FEN[3160]), .op(N5194_t0) );
fim FAN_N5194_1 ( .fault(fault), .net(N5194), .FEN(FEN[3161]), .op(N5194_t1) );
fim FAN_N5200_0 ( .fault(fault), .net(N5200), .FEN(FEN[3162]), .op(N5200_t0) );
fim FAN_N5200_1 ( .fault(fault), .net(N5200), .FEN(FEN[3163]), .op(N5200_t1) );
fim FAN_N5200_2 ( .fault(fault), .net(N5200), .FEN(FEN[3164]), .op(N5200_t2) );
fim FAN_N5206_0 ( .fault(fault), .net(N5206), .FEN(FEN[3165]), .op(N5206_t0) );
fim FAN_N5206_1 ( .fault(fault), .net(N5206), .FEN(FEN[3166]), .op(N5206_t1) );
fim FAN_N918_0 ( .fault(fault), .net(N918), .FEN(FEN[3167]), .op(N918_t0) );
fim FAN_N918_1 ( .fault(fault), .net(N918), .FEN(FEN[3168]), .op(N918_t1) );
fim FAN_N5209_0 ( .fault(fault), .net(N5209), .FEN(FEN[3169]), .op(N5209_t0) );
fim FAN_N5209_1 ( .fault(fault), .net(N5209), .FEN(FEN[3170]), .op(N5209_t1) );
fim FAN_N5209_2 ( .fault(fault), .net(N5209), .FEN(FEN[3171]), .op(N5209_t2) );
fim FAN_N5218_0 ( .fault(fault), .net(N5218), .FEN(FEN[3172]), .op(N5218_t0) );
fim FAN_N5218_1 ( .fault(fault), .net(N5218), .FEN(FEN[3173]), .op(N5218_t1) );
fim FAN_N5215_0 ( .fault(fault), .net(N5215), .FEN(FEN[3174]), .op(N5215_t0) );
fim FAN_N5215_1 ( .fault(fault), .net(N5215), .FEN(FEN[3175]), .op(N5215_t1) );
fim FAN_N5221_0 ( .fault(fault), .net(N5221), .FEN(FEN[3176]), .op(N5221_t0) );
fim FAN_N5221_1 ( .fault(fault), .net(N5221), .FEN(FEN[3177]), .op(N5221_t1) );
fim FAN_N5221_2 ( .fault(fault), .net(N5221), .FEN(FEN[3178]), .op(N5221_t2) );
fim FAN_N5227_0 ( .fault(fault), .net(N5227), .FEN(FEN[3179]), .op(N5227_t0) );
fim FAN_N5227_1 ( .fault(fault), .net(N5227), .FEN(FEN[3180]), .op(N5227_t1) );
fim FAN_N1161_0 ( .fault(fault), .net(N1161), .FEN(FEN[3181]), .op(N1161_t0) );
fim FAN_N1161_1 ( .fault(fault), .net(N1161), .FEN(FEN[3182]), .op(N1161_t1) );
fim FAN_N5230_0 ( .fault(fault), .net(N5230), .FEN(FEN[3183]), .op(N5230_t0) );
fim FAN_N5230_1 ( .fault(fault), .net(N5230), .FEN(FEN[3184]), .op(N5230_t1) );
fim FAN_N5230_2 ( .fault(fault), .net(N5230), .FEN(FEN[3185]), .op(N5230_t2) );
fim FAN_N1305_0 ( .fault(fault), .net(N1305), .FEN(FEN[3186]), .op(N1305_t0) );
fim FAN_N1305_1 ( .fault(fault), .net(N1305), .FEN(FEN[3187]), .op(N1305_t1) );
fim FAN_N5236_0 ( .fault(fault), .net(N5236), .FEN(FEN[3188]), .op(N5236_t0) );
fim FAN_N5236_1 ( .fault(fault), .net(N5236), .FEN(FEN[3189]), .op(N5236_t1) );
fim FAN_N5259_0 ( .fault(fault), .net(N5259), .FEN(FEN[3190]), .op(N5259_t0) );
fim FAN_N5259_1 ( .fault(fault), .net(N5259), .FEN(FEN[3191]), .op(N5259_t1) );
fim FAN_N5256_0 ( .fault(fault), .net(N5256), .FEN(FEN[3192]), .op(N5256_t0) );
fim FAN_N5256_1 ( .fault(fault), .net(N5256), .FEN(FEN[3193]), .op(N5256_t1) );
fim FAN_N5262_0 ( .fault(fault), .net(N5262), .FEN(FEN[3194]), .op(N5262_t0) );
fim FAN_N5262_1 ( .fault(fault), .net(N5262), .FEN(FEN[3195]), .op(N5262_t1) );
fim FAN_N5262_2 ( .fault(fault), .net(N5262), .FEN(FEN[3196]), .op(N5262_t2) );
fim FAN_N5268_0 ( .fault(fault), .net(N5268), .FEN(FEN[3197]), .op(N5268_t0) );
fim FAN_N5268_1 ( .fault(fault), .net(N5268), .FEN(FEN[3198]), .op(N5268_t1) );
fim FAN_N870_0 ( .fault(fault), .net(N870), .FEN(FEN[3199]), .op(N870_t0) );
fim FAN_N870_1 ( .fault(fault), .net(N870), .FEN(FEN[3200]), .op(N870_t1) );
fim FAN_N5271_0 ( .fault(fault), .net(N5271), .FEN(FEN[3201]), .op(N5271_t0) );
fim FAN_N5271_1 ( .fault(fault), .net(N5271), .FEN(FEN[3202]), .op(N5271_t1) );
fim FAN_N5271_2 ( .fault(fault), .net(N5271), .FEN(FEN[3203]), .op(N5271_t2) );
fim FAN_N5280_0 ( .fault(fault), .net(N5280), .FEN(FEN[3204]), .op(N5280_t0) );
fim FAN_N5280_1 ( .fault(fault), .net(N5280), .FEN(FEN[3205]), .op(N5280_t1) );
fim FAN_N5277_0 ( .fault(fault), .net(N5277), .FEN(FEN[3206]), .op(N5277_t0) );
fim FAN_N5277_1 ( .fault(fault), .net(N5277), .FEN(FEN[3207]), .op(N5277_t1) );
fim FAN_N5283_0 ( .fault(fault), .net(N5283), .FEN(FEN[3208]), .op(N5283_t0) );
fim FAN_N5283_1 ( .fault(fault), .net(N5283), .FEN(FEN[3209]), .op(N5283_t1) );
fim FAN_N5283_2 ( .fault(fault), .net(N5283), .FEN(FEN[3210]), .op(N5283_t2) );
fim FAN_N5289_0 ( .fault(fault), .net(N5289), .FEN(FEN[3211]), .op(N5289_t0) );
fim FAN_N5289_1 ( .fault(fault), .net(N5289), .FEN(FEN[3212]), .op(N5289_t1) );
fim FAN_N1113_0 ( .fault(fault), .net(N1113), .FEN(FEN[3213]), .op(N1113_t0) );
fim FAN_N1113_1 ( .fault(fault), .net(N1113), .FEN(FEN[3214]), .op(N1113_t1) );
fim FAN_N5292_0 ( .fault(fault), .net(N5292), .FEN(FEN[3215]), .op(N5292_t0) );
fim FAN_N5292_1 ( .fault(fault), .net(N5292), .FEN(FEN[3216]), .op(N5292_t1) );
fim FAN_N5292_2 ( .fault(fault), .net(N5292), .FEN(FEN[3217]), .op(N5292_t2) );
fim FAN_N5301_0 ( .fault(fault), .net(N5301), .FEN(FEN[3218]), .op(N5301_t0) );
fim FAN_N5301_1 ( .fault(fault), .net(N5301), .FEN(FEN[3219]), .op(N5301_t1) );
fim FAN_N5298_0 ( .fault(fault), .net(N5298), .FEN(FEN[3220]), .op(N5298_t0) );
fim FAN_N5298_1 ( .fault(fault), .net(N5298), .FEN(FEN[3221]), .op(N5298_t1) );
fim FAN_N5304_0 ( .fault(fault), .net(N5304), .FEN(FEN[3222]), .op(N5304_t0) );
fim FAN_N5304_1 ( .fault(fault), .net(N5304), .FEN(FEN[3223]), .op(N5304_t1) );
fim FAN_N5304_2 ( .fault(fault), .net(N5304), .FEN(FEN[3224]), .op(N5304_t2) );
fim FAN_N5309_0 ( .fault(fault), .net(N5309), .FEN(FEN[3225]), .op(N5309_t0) );
fim FAN_N5309_1 ( .fault(fault), .net(N5309), .FEN(FEN[3226]), .op(N5309_t1) );
fim FAN_N5241_0 ( .fault(fault), .net(N5241), .FEN(FEN[3227]), .op(N5241_t0) );
fim FAN_N5241_1 ( .fault(fault), .net(N5241), .FEN(FEN[3228]), .op(N5241_t1) );
fim FAN_N5312_0 ( .fault(fault), .net(N5312), .FEN(FEN[3229]), .op(N5312_t0) );
fim FAN_N5312_1 ( .fault(fault), .net(N5312), .FEN(FEN[3230]), .op(N5312_t1) );
fim FAN_N5246_0 ( .fault(fault), .net(N5246), .FEN(FEN[3231]), .op(N5246_t0) );
fim FAN_N5246_1 ( .fault(fault), .net(N5246), .FEN(FEN[3232]), .op(N5246_t1) );
fim FAN_N5315_0 ( .fault(fault), .net(N5315), .FEN(FEN[3233]), .op(N5315_t0) );
fim FAN_N5315_1 ( .fault(fault), .net(N5315), .FEN(FEN[3234]), .op(N5315_t1) );
fim FAN_N5251_0 ( .fault(fault), .net(N5251), .FEN(FEN[3235]), .op(N5251_t0) );
fim FAN_N5251_1 ( .fault(fault), .net(N5251), .FEN(FEN[3236]), .op(N5251_t1) );
fim FAN_N5318_0 ( .fault(fault), .net(N5318), .FEN(FEN[3237]), .op(N5318_t0) );
fim FAN_N5318_1 ( .fault(fault), .net(N5318), .FEN(FEN[3238]), .op(N5318_t1) );
fim FAN_N5318_2 ( .fault(fault), .net(N5318), .FEN(FEN[3239]), .op(N5318_t2) );
fim FAN_N5324_0 ( .fault(fault), .net(N5324), .FEN(FEN[3240]), .op(N5324_t0) );
fim FAN_N5324_1 ( .fault(fault), .net(N5324), .FEN(FEN[3241]), .op(N5324_t1) );
fim FAN_N822_0 ( .fault(fault), .net(N822), .FEN(FEN[3242]), .op(N822_t0) );
fim FAN_N822_1 ( .fault(fault), .net(N822), .FEN(FEN[3243]), .op(N822_t1) );
fim FAN_N5327_0 ( .fault(fault), .net(N5327), .FEN(FEN[3244]), .op(N5327_t0) );
fim FAN_N5327_1 ( .fault(fault), .net(N5327), .FEN(FEN[3245]), .op(N5327_t1) );
fim FAN_N5327_2 ( .fault(fault), .net(N5327), .FEN(FEN[3246]), .op(N5327_t2) );
fim FAN_N5336_0 ( .fault(fault), .net(N5336), .FEN(FEN[3247]), .op(N5336_t0) );
fim FAN_N5336_1 ( .fault(fault), .net(N5336), .FEN(FEN[3248]), .op(N5336_t1) );
fim FAN_N5333_0 ( .fault(fault), .net(N5333), .FEN(FEN[3249]), .op(N5333_t0) );
fim FAN_N5333_1 ( .fault(fault), .net(N5333), .FEN(FEN[3250]), .op(N5333_t1) );
fim FAN_N5339_0 ( .fault(fault), .net(N5339), .FEN(FEN[3251]), .op(N5339_t0) );
fim FAN_N5339_1 ( .fault(fault), .net(N5339), .FEN(FEN[3252]), .op(N5339_t1) );
fim FAN_N5339_2 ( .fault(fault), .net(N5339), .FEN(FEN[3253]), .op(N5339_t2) );
fim FAN_N5345_0 ( .fault(fault), .net(N5345), .FEN(FEN[3254]), .op(N5345_t0) );
fim FAN_N5345_1 ( .fault(fault), .net(N5345), .FEN(FEN[3255]), .op(N5345_t1) );
fim FAN_N1065_0 ( .fault(fault), .net(N1065), .FEN(FEN[3256]), .op(N1065_t0) );
fim FAN_N1065_1 ( .fault(fault), .net(N1065), .FEN(FEN[3257]), .op(N1065_t1) );
fim FAN_N5348_0 ( .fault(fault), .net(N5348), .FEN(FEN[3258]), .op(N5348_t0) );
fim FAN_N5348_1 ( .fault(fault), .net(N5348), .FEN(FEN[3259]), .op(N5348_t1) );
fim FAN_N5348_2 ( .fault(fault), .net(N5348), .FEN(FEN[3260]), .op(N5348_t2) );
fim FAN_N5357_0 ( .fault(fault), .net(N5357), .FEN(FEN[3261]), .op(N5357_t0) );
fim FAN_N5357_1 ( .fault(fault), .net(N5357), .FEN(FEN[3262]), .op(N5357_t1) );
fim FAN_N5354_0 ( .fault(fault), .net(N5354), .FEN(FEN[3263]), .op(N5354_t0) );
fim FAN_N5354_1 ( .fault(fault), .net(N5354), .FEN(FEN[3264]), .op(N5354_t1) );
fim FAN_N5360_0 ( .fault(fault), .net(N5360), .FEN(FEN[3265]), .op(N5360_t0) );
fim FAN_N5360_1 ( .fault(fault), .net(N5360), .FEN(FEN[3266]), .op(N5360_t1) );
fim FAN_N5360_2 ( .fault(fault), .net(N5360), .FEN(FEN[3267]), .op(N5360_t2) );
fim FAN_N5366_0 ( .fault(fault), .net(N5366), .FEN(FEN[3268]), .op(N5366_t0) );
fim FAN_N5366_1 ( .fault(fault), .net(N5366), .FEN(FEN[3269]), .op(N5366_t1) );
fim FAN_N5366_2 ( .fault(fault), .net(N5366), .FEN(FEN[3270]), .op(N5366_t2) );
fim FAN_N5370_0 ( .fault(fault), .net(N5370), .FEN(FEN[3271]), .op(N5370_t0) );
fim FAN_N5370_1 ( .fault(fault), .net(N5370), .FEN(FEN[3272]), .op(N5370_t1) );
fim FAN_N5370_2 ( .fault(fault), .net(N5370), .FEN(FEN[3273]), .op(N5370_t2) );
fim FAN_N5374_0 ( .fault(fault), .net(N5374), .FEN(FEN[3274]), .op(N5374_t0) );
fim FAN_N5374_1 ( .fault(fault), .net(N5374), .FEN(FEN[3275]), .op(N5374_t1) );
fim FAN_N5374_2 ( .fault(fault), .net(N5374), .FEN(FEN[3276]), .op(N5374_t2) );
fim FAN_N5380_0 ( .fault(fault), .net(N5380), .FEN(FEN[3277]), .op(N5380_t0) );
fim FAN_N5380_1 ( .fault(fault), .net(N5380), .FEN(FEN[3278]), .op(N5380_t1) );
fim FAN_N774_0 ( .fault(fault), .net(N774), .FEN(FEN[3279]), .op(N774_t0) );
fim FAN_N774_1 ( .fault(fault), .net(N774), .FEN(FEN[3280]), .op(N774_t1) );
fim FAN_N5383_0 ( .fault(fault), .net(N5383), .FEN(FEN[3281]), .op(N5383_t0) );
fim FAN_N5383_1 ( .fault(fault), .net(N5383), .FEN(FEN[3282]), .op(N5383_t1) );
fim FAN_N5383_2 ( .fault(fault), .net(N5383), .FEN(FEN[3283]), .op(N5383_t2) );
fim FAN_N5392_0 ( .fault(fault), .net(N5392), .FEN(FEN[3284]), .op(N5392_t0) );
fim FAN_N5392_1 ( .fault(fault), .net(N5392), .FEN(FEN[3285]), .op(N5392_t1) );
fim FAN_N5389_0 ( .fault(fault), .net(N5389), .FEN(FEN[3286]), .op(N5389_t0) );
fim FAN_N5389_1 ( .fault(fault), .net(N5389), .FEN(FEN[3287]), .op(N5389_t1) );
fim FAN_N5395_0 ( .fault(fault), .net(N5395), .FEN(FEN[3288]), .op(N5395_t0) );
fim FAN_N5395_1 ( .fault(fault), .net(N5395), .FEN(FEN[3289]), .op(N5395_t1) );
fim FAN_N5395_2 ( .fault(fault), .net(N5395), .FEN(FEN[3290]), .op(N5395_t2) );
fim FAN_N5401_0 ( .fault(fault), .net(N5401), .FEN(FEN[3291]), .op(N5401_t0) );
fim FAN_N5401_1 ( .fault(fault), .net(N5401), .FEN(FEN[3292]), .op(N5401_t1) );
fim FAN_N1017_0 ( .fault(fault), .net(N1017), .FEN(FEN[3293]), .op(N1017_t0) );
fim FAN_N1017_1 ( .fault(fault), .net(N1017), .FEN(FEN[3294]), .op(N1017_t1) );
fim FAN_N5404_0 ( .fault(fault), .net(N5404), .FEN(FEN[3295]), .op(N5404_t0) );
fim FAN_N5404_1 ( .fault(fault), .net(N5404), .FEN(FEN[3296]), .op(N5404_t1) );
fim FAN_N5404_2 ( .fault(fault), .net(N5404), .FEN(FEN[3297]), .op(N5404_t2) );
fim FAN_N5413_0 ( .fault(fault), .net(N5413), .FEN(FEN[3298]), .op(N5413_t0) );
fim FAN_N5413_1 ( .fault(fault), .net(N5413), .FEN(FEN[3299]), .op(N5413_t1) );
fim FAN_N5410_0 ( .fault(fault), .net(N5410), .FEN(FEN[3300]), .op(N5410_t0) );
fim FAN_N5410_1 ( .fault(fault), .net(N5410), .FEN(FEN[3301]), .op(N5410_t1) );
fim FAN_N5416_0 ( .fault(fault), .net(N5416), .FEN(FEN[3302]), .op(N5416_t0) );
fim FAN_N5416_1 ( .fault(fault), .net(N5416), .FEN(FEN[3303]), .op(N5416_t1) );
fim FAN_N5416_2 ( .fault(fault), .net(N5416), .FEN(FEN[3304]), .op(N5416_t2) );
fim FAN_N5422_0 ( .fault(fault), .net(N5422), .FEN(FEN[3305]), .op(N5422_t0) );
fim FAN_N5422_1 ( .fault(fault), .net(N5422), .FEN(FEN[3306]), .op(N5422_t1) );
fim FAN_N1260_0 ( .fault(fault), .net(N1260), .FEN(FEN[3307]), .op(N1260_t0) );
fim FAN_N1260_1 ( .fault(fault), .net(N1260), .FEN(FEN[3308]), .op(N1260_t1) );
fim FAN_N5431_0 ( .fault(fault), .net(N5431), .FEN(FEN[3309]), .op(N5431_t0) );
fim FAN_N5431_1 ( .fault(fault), .net(N5431), .FEN(FEN[3310]), .op(N5431_t1) );
fim FAN_N726_0 ( .fault(fault), .net(N726), .FEN(FEN[3311]), .op(N726_t0) );
fim FAN_N726_1 ( .fault(fault), .net(N726), .FEN(FEN[3312]), .op(N726_t1) );
fim FAN_N5434_0 ( .fault(fault), .net(N5434), .FEN(FEN[3313]), .op(N5434_t0) );
fim FAN_N5434_1 ( .fault(fault), .net(N5434), .FEN(FEN[3314]), .op(N5434_t1) );
fim FAN_N5434_2 ( .fault(fault), .net(N5434), .FEN(FEN[3315]), .op(N5434_t2) );
fim FAN_N5443_0 ( .fault(fault), .net(N5443), .FEN(FEN[3316]), .op(N5443_t0) );
fim FAN_N5443_1 ( .fault(fault), .net(N5443), .FEN(FEN[3317]), .op(N5443_t1) );
fim FAN_N5440_0 ( .fault(fault), .net(N5440), .FEN(FEN[3318]), .op(N5440_t0) );
fim FAN_N5440_1 ( .fault(fault), .net(N5440), .FEN(FEN[3319]), .op(N5440_t1) );
fim FAN_N5446_0 ( .fault(fault), .net(N5446), .FEN(FEN[3320]), .op(N5446_t0) );
fim FAN_N5446_1 ( .fault(fault), .net(N5446), .FEN(FEN[3321]), .op(N5446_t1) );
fim FAN_N5446_2 ( .fault(fault), .net(N5446), .FEN(FEN[3322]), .op(N5446_t2) );
fim FAN_N5452_0 ( .fault(fault), .net(N5452), .FEN(FEN[3323]), .op(N5452_t0) );
fim FAN_N5452_1 ( .fault(fault), .net(N5452), .FEN(FEN[3324]), .op(N5452_t1) );
fim FAN_N969_0 ( .fault(fault), .net(N969), .FEN(FEN[3325]), .op(N969_t0) );
fim FAN_N969_1 ( .fault(fault), .net(N969), .FEN(FEN[3326]), .op(N969_t1) );
fim FAN_N5455_0 ( .fault(fault), .net(N5455), .FEN(FEN[3327]), .op(N5455_t0) );
fim FAN_N5455_1 ( .fault(fault), .net(N5455), .FEN(FEN[3328]), .op(N5455_t1) );
fim FAN_N5455_2 ( .fault(fault), .net(N5455), .FEN(FEN[3329]), .op(N5455_t2) );
fim FAN_N5464_0 ( .fault(fault), .net(N5464), .FEN(FEN[3330]), .op(N5464_t0) );
fim FAN_N5464_1 ( .fault(fault), .net(N5464), .FEN(FEN[3331]), .op(N5464_t1) );
fim FAN_N5461_0 ( .fault(fault), .net(N5461), .FEN(FEN[3332]), .op(N5461_t0) );
fim FAN_N5461_1 ( .fault(fault), .net(N5461), .FEN(FEN[3333]), .op(N5461_t1) );
fim FAN_N5467_0 ( .fault(fault), .net(N5467), .FEN(FEN[3334]), .op(N5467_t0) );
fim FAN_N5467_1 ( .fault(fault), .net(N5467), .FEN(FEN[3335]), .op(N5467_t1) );
fim FAN_N5467_2 ( .fault(fault), .net(N5467), .FEN(FEN[3336]), .op(N5467_t2) );
fim FAN_N5473_0 ( .fault(fault), .net(N5473), .FEN(FEN[3337]), .op(N5473_t0) );
fim FAN_N5473_1 ( .fault(fault), .net(N5473), .FEN(FEN[3338]), .op(N5473_t1) );
fim FAN_N1212_0 ( .fault(fault), .net(N1212), .FEN(FEN[3339]), .op(N1212_t0) );
fim FAN_N1212_1 ( .fault(fault), .net(N1212), .FEN(FEN[3340]), .op(N1212_t1) );
fim FAN_N5476_0 ( .fault(fault), .net(N5476), .FEN(FEN[3341]), .op(N5476_t0) );
fim FAN_N5476_1 ( .fault(fault), .net(N5476), .FEN(FEN[3342]), .op(N5476_t1) );
fim FAN_N5476_2 ( .fault(fault), .net(N5476), .FEN(FEN[3343]), .op(N5476_t2) );
fim FAN_N5480_0 ( .fault(fault), .net(N5480), .FEN(FEN[3344]), .op(N5480_t0) );
fim FAN_N5480_1 ( .fault(fault), .net(N5480), .FEN(FEN[3345]), .op(N5480_t1) );
fim FAN_N582_0 ( .fault(fault), .net(N582), .FEN(FEN[3346]), .op(N582_t0) );
fim FAN_N582_1 ( .fault(fault), .net(N582), .FEN(FEN[3347]), .op(N582_t1) );
fim FAN_N5483_0 ( .fault(fault), .net(N5483), .FEN(FEN[3348]), .op(N5483_t0) );
fim FAN_N5483_1 ( .fault(fault), .net(N5483), .FEN(FEN[3349]), .op(N5483_t1) );
fim FAN_N630_0 ( .fault(fault), .net(N630), .FEN(FEN[3350]), .op(N630_t0) );
fim FAN_N630_1 ( .fault(fault), .net(N630), .FEN(FEN[3351]), .op(N630_t1) );
fim FAN_N5486_0 ( .fault(fault), .net(N5486), .FEN(FEN[3352]), .op(N5486_t0) );
fim FAN_N5486_1 ( .fault(fault), .net(N5486), .FEN(FEN[3353]), .op(N5486_t1) );
fim FAN_N678_0 ( .fault(fault), .net(N678), .FEN(FEN[3354]), .op(N678_t0) );
fim FAN_N678_1 ( .fault(fault), .net(N678), .FEN(FEN[3355]), .op(N678_t1) );
fim FAN_N5489_0 ( .fault(fault), .net(N5489), .FEN(FEN[3356]), .op(N5489_t0) );
fim FAN_N5489_1 ( .fault(fault), .net(N5489), .FEN(FEN[3357]), .op(N5489_t1) );
fim FAN_N5489_2 ( .fault(fault), .net(N5489), .FEN(FEN[3358]), .op(N5489_t2) );
fim FAN_N5498_0 ( .fault(fault), .net(N5498), .FEN(FEN[3359]), .op(N5498_t0) );
fim FAN_N5498_1 ( .fault(fault), .net(N5498), .FEN(FEN[3360]), .op(N5498_t1) );
fim FAN_N5495_0 ( .fault(fault), .net(N5495), .FEN(FEN[3361]), .op(N5495_t0) );
fim FAN_N5495_1 ( .fault(fault), .net(N5495), .FEN(FEN[3362]), .op(N5495_t1) );
fim FAN_N5501_0 ( .fault(fault), .net(N5501), .FEN(FEN[3363]), .op(N5501_t0) );
fim FAN_N5501_1 ( .fault(fault), .net(N5501), .FEN(FEN[3364]), .op(N5501_t1) );
fim FAN_N5501_2 ( .fault(fault), .net(N5501), .FEN(FEN[3365]), .op(N5501_t2) );
fim FAN_N5507_0 ( .fault(fault), .net(N5507), .FEN(FEN[3366]), .op(N5507_t0) );
fim FAN_N5507_1 ( .fault(fault), .net(N5507), .FEN(FEN[3367]), .op(N5507_t1) );
fim FAN_N921_0 ( .fault(fault), .net(N921), .FEN(FEN[3368]), .op(N921_t0) );
fim FAN_N921_1 ( .fault(fault), .net(N921), .FEN(FEN[3369]), .op(N921_t1) );
fim FAN_N5510_0 ( .fault(fault), .net(N5510), .FEN(FEN[3370]), .op(N5510_t0) );
fim FAN_N5510_1 ( .fault(fault), .net(N5510), .FEN(FEN[3371]), .op(N5510_t1) );
fim FAN_N5510_2 ( .fault(fault), .net(N5510), .FEN(FEN[3372]), .op(N5510_t2) );
fim FAN_N5519_0 ( .fault(fault), .net(N5519), .FEN(FEN[3373]), .op(N5519_t0) );
fim FAN_N5519_1 ( .fault(fault), .net(N5519), .FEN(FEN[3374]), .op(N5519_t1) );
fim FAN_N5516_0 ( .fault(fault), .net(N5516), .FEN(FEN[3375]), .op(N5516_t0) );
fim FAN_N5516_1 ( .fault(fault), .net(N5516), .FEN(FEN[3376]), .op(N5516_t1) );
fim FAN_N5522_0 ( .fault(fault), .net(N5522), .FEN(FEN[3377]), .op(N5522_t0) );
fim FAN_N5522_1 ( .fault(fault), .net(N5522), .FEN(FEN[3378]), .op(N5522_t1) );
fim FAN_N5522_2 ( .fault(fault), .net(N5522), .FEN(FEN[3379]), .op(N5522_t2) );
fim FAN_N5528_0 ( .fault(fault), .net(N5528), .FEN(FEN[3380]), .op(N5528_t0) );
fim FAN_N5528_1 ( .fault(fault), .net(N5528), .FEN(FEN[3381]), .op(N5528_t1) );
fim FAN_N1164_0 ( .fault(fault), .net(N1164), .FEN(FEN[3382]), .op(N1164_t0) );
fim FAN_N1164_1 ( .fault(fault), .net(N1164), .FEN(FEN[3383]), .op(N1164_t1) );
fim FAN_N5531_0 ( .fault(fault), .net(N5531), .FEN(FEN[3384]), .op(N5531_t0) );
fim FAN_N5531_1 ( .fault(fault), .net(N5531), .FEN(FEN[3385]), .op(N5531_t1) );
fim FAN_N5531_2 ( .fault(fault), .net(N5531), .FEN(FEN[3386]), .op(N5531_t2) );
fim FAN_N1308_0 ( .fault(fault), .net(N1308), .FEN(FEN[3387]), .op(N1308_t0) );
fim FAN_N1308_1 ( .fault(fault), .net(N1308), .FEN(FEN[3388]), .op(N1308_t1) );
fim FAN_N5537_0 ( .fault(fault), .net(N5537), .FEN(FEN[3389]), .op(N5537_t0) );
fim FAN_N5537_1 ( .fault(fault), .net(N5537), .FEN(FEN[3390]), .op(N5537_t1) );
fim FAN_N5540_0 ( .fault(fault), .net(N5540), .FEN(FEN[3391]), .op(N5540_t0) );
fim FAN_N5540_1 ( .fault(fault), .net(N5540), .FEN(FEN[3392]), .op(N5540_t1) );
fim FAN_N5540_2 ( .fault(fault), .net(N5540), .FEN(FEN[3393]), .op(N5540_t2) );
fim FAN_N5544_0 ( .fault(fault), .net(N5544), .FEN(FEN[3394]), .op(N5544_t0) );
fim FAN_N5544_1 ( .fault(fault), .net(N5544), .FEN(FEN[3395]), .op(N5544_t1) );
fim FAN_N5544_2 ( .fault(fault), .net(N5544), .FEN(FEN[3396]), .op(N5544_t2) );
fim FAN_N5548_0 ( .fault(fault), .net(N5548), .FEN(FEN[3397]), .op(N5548_t0) );
fim FAN_N5548_1 ( .fault(fault), .net(N5548), .FEN(FEN[3398]), .op(N5548_t1) );
fim FAN_N5548_2 ( .fault(fault), .net(N5548), .FEN(FEN[3399]), .op(N5548_t2) );
fim FAN_N5557_0 ( .fault(fault), .net(N5557), .FEN(FEN[3400]), .op(N5557_t0) );
fim FAN_N5557_1 ( .fault(fault), .net(N5557), .FEN(FEN[3401]), .op(N5557_t1) );
fim FAN_N5554_0 ( .fault(fault), .net(N5554), .FEN(FEN[3402]), .op(N5554_t0) );
fim FAN_N5554_1 ( .fault(fault), .net(N5554), .FEN(FEN[3403]), .op(N5554_t1) );
fim FAN_N5560_0 ( .fault(fault), .net(N5560), .FEN(FEN[3404]), .op(N5560_t0) );
fim FAN_N5560_1 ( .fault(fault), .net(N5560), .FEN(FEN[3405]), .op(N5560_t1) );
fim FAN_N5560_2 ( .fault(fault), .net(N5560), .FEN(FEN[3406]), .op(N5560_t2) );
fim FAN_N5566_0 ( .fault(fault), .net(N5566), .FEN(FEN[3407]), .op(N5566_t0) );
fim FAN_N5566_1 ( .fault(fault), .net(N5566), .FEN(FEN[3408]), .op(N5566_t1) );
fim FAN_N873_0 ( .fault(fault), .net(N873), .FEN(FEN[3409]), .op(N873_t0) );
fim FAN_N873_1 ( .fault(fault), .net(N873), .FEN(FEN[3410]), .op(N873_t1) );
fim FAN_N5569_0 ( .fault(fault), .net(N5569), .FEN(FEN[3411]), .op(N5569_t0) );
fim FAN_N5569_1 ( .fault(fault), .net(N5569), .FEN(FEN[3412]), .op(N5569_t1) );
fim FAN_N5569_2 ( .fault(fault), .net(N5569), .FEN(FEN[3413]), .op(N5569_t2) );
fim FAN_N5578_0 ( .fault(fault), .net(N5578), .FEN(FEN[3414]), .op(N5578_t0) );
fim FAN_N5578_1 ( .fault(fault), .net(N5578), .FEN(FEN[3415]), .op(N5578_t1) );
fim FAN_N5575_0 ( .fault(fault), .net(N5575), .FEN(FEN[3416]), .op(N5575_t0) );
fim FAN_N5575_1 ( .fault(fault), .net(N5575), .FEN(FEN[3417]), .op(N5575_t1) );
fim FAN_N5581_0 ( .fault(fault), .net(N5581), .FEN(FEN[3418]), .op(N5581_t0) );
fim FAN_N5581_1 ( .fault(fault), .net(N5581), .FEN(FEN[3419]), .op(N5581_t1) );
fim FAN_N5581_2 ( .fault(fault), .net(N5581), .FEN(FEN[3420]), .op(N5581_t2) );
fim FAN_N5587_0 ( .fault(fault), .net(N5587), .FEN(FEN[3421]), .op(N5587_t0) );
fim FAN_N5587_1 ( .fault(fault), .net(N5587), .FEN(FEN[3422]), .op(N5587_t1) );
fim FAN_N1116_0 ( .fault(fault), .net(N1116), .FEN(FEN[3423]), .op(N1116_t0) );
fim FAN_N1116_1 ( .fault(fault), .net(N1116), .FEN(FEN[3424]), .op(N1116_t1) );
fim FAN_N5590_0 ( .fault(fault), .net(N5590), .FEN(FEN[3425]), .op(N5590_t0) );
fim FAN_N5590_1 ( .fault(fault), .net(N5590), .FEN(FEN[3426]), .op(N5590_t1) );
fim FAN_N5590_2 ( .fault(fault), .net(N5590), .FEN(FEN[3427]), .op(N5590_t2) );
fim FAN_N5599_0 ( .fault(fault), .net(N5599), .FEN(FEN[3428]), .op(N5599_t0) );
fim FAN_N5599_1 ( .fault(fault), .net(N5599), .FEN(FEN[3429]), .op(N5599_t1) );
fim FAN_N5596_0 ( .fault(fault), .net(N5596), .FEN(FEN[3430]), .op(N5596_t0) );
fim FAN_N5596_1 ( .fault(fault), .net(N5596), .FEN(FEN[3431]), .op(N5596_t1) );
fim FAN_N5602_0 ( .fault(fault), .net(N5602), .FEN(FEN[3432]), .op(N5602_t0) );
fim FAN_N5602_1 ( .fault(fault), .net(N5602), .FEN(FEN[3433]), .op(N5602_t1) );
fim FAN_N5602_2 ( .fault(fault), .net(N5602), .FEN(FEN[3434]), .op(N5602_t2) );
fim FAN_N5621_0 ( .fault(fault), .net(N5621), .FEN(FEN[3435]), .op(N5621_t0) );
fim FAN_N5621_1 ( .fault(fault), .net(N5621), .FEN(FEN[3436]), .op(N5621_t1) );
fim FAN_N5618_0 ( .fault(fault), .net(N5618), .FEN(FEN[3437]), .op(N5618_t0) );
fim FAN_N5618_1 ( .fault(fault), .net(N5618), .FEN(FEN[3438]), .op(N5618_t1) );
fim FAN_N5624_0 ( .fault(fault), .net(N5624), .FEN(FEN[3439]), .op(N5624_t0) );
fim FAN_N5624_1 ( .fault(fault), .net(N5624), .FEN(FEN[3440]), .op(N5624_t1) );
fim FAN_N5624_2 ( .fault(fault), .net(N5624), .FEN(FEN[3441]), .op(N5624_t2) );
fim FAN_N5630_0 ( .fault(fault), .net(N5630), .FEN(FEN[3442]), .op(N5630_t0) );
fim FAN_N5630_1 ( .fault(fault), .net(N5630), .FEN(FEN[3443]), .op(N5630_t1) );
fim FAN_N825_0 ( .fault(fault), .net(N825), .FEN(FEN[3444]), .op(N825_t0) );
fim FAN_N825_1 ( .fault(fault), .net(N825), .FEN(FEN[3445]), .op(N825_t1) );
fim FAN_N5633_0 ( .fault(fault), .net(N5633), .FEN(FEN[3446]), .op(N5633_t0) );
fim FAN_N5633_1 ( .fault(fault), .net(N5633), .FEN(FEN[3447]), .op(N5633_t1) );
fim FAN_N5633_2 ( .fault(fault), .net(N5633), .FEN(FEN[3448]), .op(N5633_t2) );
fim FAN_N5642_0 ( .fault(fault), .net(N5642), .FEN(FEN[3449]), .op(N5642_t0) );
fim FAN_N5642_1 ( .fault(fault), .net(N5642), .FEN(FEN[3450]), .op(N5642_t1) );
fim FAN_N5639_0 ( .fault(fault), .net(N5639), .FEN(FEN[3451]), .op(N5639_t0) );
fim FAN_N5639_1 ( .fault(fault), .net(N5639), .FEN(FEN[3452]), .op(N5639_t1) );
fim FAN_N5645_0 ( .fault(fault), .net(N5645), .FEN(FEN[3453]), .op(N5645_t0) );
fim FAN_N5645_1 ( .fault(fault), .net(N5645), .FEN(FEN[3454]), .op(N5645_t1) );
fim FAN_N5645_2 ( .fault(fault), .net(N5645), .FEN(FEN[3455]), .op(N5645_t2) );
fim FAN_N5651_0 ( .fault(fault), .net(N5651), .FEN(FEN[3456]), .op(N5651_t0) );
fim FAN_N5651_1 ( .fault(fault), .net(N5651), .FEN(FEN[3457]), .op(N5651_t1) );
fim FAN_N1068_0 ( .fault(fault), .net(N1068), .FEN(FEN[3458]), .op(N1068_t0) );
fim FAN_N1068_1 ( .fault(fault), .net(N1068), .FEN(FEN[3459]), .op(N1068_t1) );
fim FAN_N5654_0 ( .fault(fault), .net(N5654), .FEN(FEN[3460]), .op(N5654_t0) );
fim FAN_N5654_1 ( .fault(fault), .net(N5654), .FEN(FEN[3461]), .op(N5654_t1) );
fim FAN_N5654_2 ( .fault(fault), .net(N5654), .FEN(FEN[3462]), .op(N5654_t2) );
fim FAN_N5663_0 ( .fault(fault), .net(N5663), .FEN(FEN[3463]), .op(N5663_t0) );
fim FAN_N5663_1 ( .fault(fault), .net(N5663), .FEN(FEN[3464]), .op(N5663_t1) );
fim FAN_N5660_0 ( .fault(fault), .net(N5660), .FEN(FEN[3465]), .op(N5660_t0) );
fim FAN_N5660_1 ( .fault(fault), .net(N5660), .FEN(FEN[3466]), .op(N5660_t1) );
fim FAN_N5666_0 ( .fault(fault), .net(N5666), .FEN(FEN[3467]), .op(N5666_t0) );
fim FAN_N5666_1 ( .fault(fault), .net(N5666), .FEN(FEN[3468]), .op(N5666_t1) );
fim FAN_N5666_2 ( .fault(fault), .net(N5666), .FEN(FEN[3469]), .op(N5666_t2) );
fim FAN_N5673_0 ( .fault(fault), .net(N5673), .FEN(FEN[3470]), .op(N5673_t0) );
fim FAN_N5673_1 ( .fault(fault), .net(N5673), .FEN(FEN[3471]), .op(N5673_t1) );
fim FAN_N5608_0 ( .fault(fault), .net(N5608), .FEN(FEN[3472]), .op(N5608_t0) );
fim FAN_N5608_1 ( .fault(fault), .net(N5608), .FEN(FEN[3473]), .op(N5608_t1) );
fim FAN_N5676_0 ( .fault(fault), .net(N5676), .FEN(FEN[3474]), .op(N5676_t0) );
fim FAN_N5676_1 ( .fault(fault), .net(N5676), .FEN(FEN[3475]), .op(N5676_t1) );
fim FAN_N5613_0 ( .fault(fault), .net(N5613), .FEN(FEN[3476]), .op(N5613_t0) );
fim FAN_N5613_1 ( .fault(fault), .net(N5613), .FEN(FEN[3477]), .op(N5613_t1) );
fim FAN_N5679_0 ( .fault(fault), .net(N5679), .FEN(FEN[3478]), .op(N5679_t0) );
fim FAN_N5679_1 ( .fault(fault), .net(N5679), .FEN(FEN[3479]), .op(N5679_t1) );
fim FAN_N5679_2 ( .fault(fault), .net(N5679), .FEN(FEN[3480]), .op(N5679_t2) );
fim FAN_N5685_0 ( .fault(fault), .net(N5685), .FEN(FEN[3481]), .op(N5685_t0) );
fim FAN_N5685_1 ( .fault(fault), .net(N5685), .FEN(FEN[3482]), .op(N5685_t1) );
fim FAN_N777_0 ( .fault(fault), .net(N777), .FEN(FEN[3483]), .op(N777_t0) );
fim FAN_N777_1 ( .fault(fault), .net(N777), .FEN(FEN[3484]), .op(N777_t1) );
fim FAN_N5688_0 ( .fault(fault), .net(N5688), .FEN(FEN[3485]), .op(N5688_t0) );
fim FAN_N5688_1 ( .fault(fault), .net(N5688), .FEN(FEN[3486]), .op(N5688_t1) );
fim FAN_N5688_2 ( .fault(fault), .net(N5688), .FEN(FEN[3487]), .op(N5688_t2) );
fim FAN_N5697_0 ( .fault(fault), .net(N5697), .FEN(FEN[3488]), .op(N5697_t0) );
fim FAN_N5697_1 ( .fault(fault), .net(N5697), .FEN(FEN[3489]), .op(N5697_t1) );
fim FAN_N5694_0 ( .fault(fault), .net(N5694), .FEN(FEN[3490]), .op(N5694_t0) );
fim FAN_N5694_1 ( .fault(fault), .net(N5694), .FEN(FEN[3491]), .op(N5694_t1) );
fim FAN_N5700_0 ( .fault(fault), .net(N5700), .FEN(FEN[3492]), .op(N5700_t0) );
fim FAN_N5700_1 ( .fault(fault), .net(N5700), .FEN(FEN[3493]), .op(N5700_t1) );
fim FAN_N5700_2 ( .fault(fault), .net(N5700), .FEN(FEN[3494]), .op(N5700_t2) );
fim FAN_N5706_0 ( .fault(fault), .net(N5706), .FEN(FEN[3495]), .op(N5706_t0) );
fim FAN_N5706_1 ( .fault(fault), .net(N5706), .FEN(FEN[3496]), .op(N5706_t1) );
fim FAN_N1020_0 ( .fault(fault), .net(N1020), .FEN(FEN[3497]), .op(N1020_t0) );
fim FAN_N1020_1 ( .fault(fault), .net(N1020), .FEN(FEN[3498]), .op(N1020_t1) );
fim FAN_N5709_0 ( .fault(fault), .net(N5709), .FEN(FEN[3499]), .op(N5709_t0) );
fim FAN_N5709_1 ( .fault(fault), .net(N5709), .FEN(FEN[3500]), .op(N5709_t1) );
fim FAN_N5709_2 ( .fault(fault), .net(N5709), .FEN(FEN[3501]), .op(N5709_t2) );
fim FAN_N5718_0 ( .fault(fault), .net(N5718), .FEN(FEN[3502]), .op(N5718_t0) );
fim FAN_N5718_1 ( .fault(fault), .net(N5718), .FEN(FEN[3503]), .op(N5718_t1) );
fim FAN_N5715_0 ( .fault(fault), .net(N5715), .FEN(FEN[3504]), .op(N5715_t0) );
fim FAN_N5715_1 ( .fault(fault), .net(N5715), .FEN(FEN[3505]), .op(N5715_t1) );
fim FAN_N5721_0 ( .fault(fault), .net(N5721), .FEN(FEN[3506]), .op(N5721_t0) );
fim FAN_N5721_1 ( .fault(fault), .net(N5721), .FEN(FEN[3507]), .op(N5721_t1) );
fim FAN_N5721_2 ( .fault(fault), .net(N5721), .FEN(FEN[3508]), .op(N5721_t2) );
fim FAN_N5730_0 ( .fault(fault), .net(N5730), .FEN(FEN[3509]), .op(N5730_t0) );
fim FAN_N5730_1 ( .fault(fault), .net(N5730), .FEN(FEN[3510]), .op(N5730_t1) );
fim FAN_N5730_2 ( .fault(fault), .net(N5730), .FEN(FEN[3511]), .op(N5730_t2) );
fim FAN_N5734_0 ( .fault(fault), .net(N5734), .FEN(FEN[3512]), .op(N5734_t0) );
fim FAN_N5734_1 ( .fault(fault), .net(N5734), .FEN(FEN[3513]), .op(N5734_t1) );
fim FAN_N5734_2 ( .fault(fault), .net(N5734), .FEN(FEN[3514]), .op(N5734_t2) );
fim FAN_N5740_0 ( .fault(fault), .net(N5740), .FEN(FEN[3515]), .op(N5740_t0) );
fim FAN_N5740_1 ( .fault(fault), .net(N5740), .FEN(FEN[3516]), .op(N5740_t1) );
fim FAN_N729_0 ( .fault(fault), .net(N729), .FEN(FEN[3517]), .op(N729_t0) );
fim FAN_N729_1 ( .fault(fault), .net(N729), .FEN(FEN[3518]), .op(N729_t1) );
fim FAN_N5743_0 ( .fault(fault), .net(N5743), .FEN(FEN[3519]), .op(N5743_t0) );
fim FAN_N5743_1 ( .fault(fault), .net(N5743), .FEN(FEN[3520]), .op(N5743_t1) );
fim FAN_N5743_2 ( .fault(fault), .net(N5743), .FEN(FEN[3521]), .op(N5743_t2) );
fim FAN_N5752_0 ( .fault(fault), .net(N5752), .FEN(FEN[3522]), .op(N5752_t0) );
fim FAN_N5752_1 ( .fault(fault), .net(N5752), .FEN(FEN[3523]), .op(N5752_t1) );
fim FAN_N5749_0 ( .fault(fault), .net(N5749), .FEN(FEN[3524]), .op(N5749_t0) );
fim FAN_N5749_1 ( .fault(fault), .net(N5749), .FEN(FEN[3525]), .op(N5749_t1) );
fim FAN_N5755_0 ( .fault(fault), .net(N5755), .FEN(FEN[3526]), .op(N5755_t0) );
fim FAN_N5755_1 ( .fault(fault), .net(N5755), .FEN(FEN[3527]), .op(N5755_t1) );
fim FAN_N5755_2 ( .fault(fault), .net(N5755), .FEN(FEN[3528]), .op(N5755_t2) );
fim FAN_N5761_0 ( .fault(fault), .net(N5761), .FEN(FEN[3529]), .op(N5761_t0) );
fim FAN_N5761_1 ( .fault(fault), .net(N5761), .FEN(FEN[3530]), .op(N5761_t1) );
fim FAN_N972_0 ( .fault(fault), .net(N972), .FEN(FEN[3531]), .op(N972_t0) );
fim FAN_N972_1 ( .fault(fault), .net(N972), .FEN(FEN[3532]), .op(N972_t1) );
fim FAN_N5764_0 ( .fault(fault), .net(N5764), .FEN(FEN[3533]), .op(N5764_t0) );
fim FAN_N5764_1 ( .fault(fault), .net(N5764), .FEN(FEN[3534]), .op(N5764_t1) );
fim FAN_N5764_2 ( .fault(fault), .net(N5764), .FEN(FEN[3535]), .op(N5764_t2) );
fim FAN_N5773_0 ( .fault(fault), .net(N5773), .FEN(FEN[3536]), .op(N5773_t0) );
fim FAN_N5773_1 ( .fault(fault), .net(N5773), .FEN(FEN[3537]), .op(N5773_t1) );
fim FAN_N5770_0 ( .fault(fault), .net(N5770), .FEN(FEN[3538]), .op(N5770_t0) );
fim FAN_N5770_1 ( .fault(fault), .net(N5770), .FEN(FEN[3539]), .op(N5770_t1) );
fim FAN_N5776_0 ( .fault(fault), .net(N5776), .FEN(FEN[3540]), .op(N5776_t0) );
fim FAN_N5776_1 ( .fault(fault), .net(N5776), .FEN(FEN[3541]), .op(N5776_t1) );
fim FAN_N5776_2 ( .fault(fault), .net(N5776), .FEN(FEN[3542]), .op(N5776_t2) );
fim FAN_N5789_0 ( .fault(fault), .net(N5789), .FEN(FEN[3543]), .op(N5789_t0) );
fim FAN_N5789_1 ( .fault(fault), .net(N5789), .FEN(FEN[3544]), .op(N5789_t1) );
fim FAN_N681_0 ( .fault(fault), .net(N681), .FEN(FEN[3545]), .op(N681_t0) );
fim FAN_N681_1 ( .fault(fault), .net(N681), .FEN(FEN[3546]), .op(N681_t1) );
fim FAN_N5792_0 ( .fault(fault), .net(N5792), .FEN(FEN[3547]), .op(N5792_t0) );
fim FAN_N5792_1 ( .fault(fault), .net(N5792), .FEN(FEN[3548]), .op(N5792_t1) );
fim FAN_N5792_2 ( .fault(fault), .net(N5792), .FEN(FEN[3549]), .op(N5792_t2) );
fim FAN_N5801_0 ( .fault(fault), .net(N5801), .FEN(FEN[3550]), .op(N5801_t0) );
fim FAN_N5801_1 ( .fault(fault), .net(N5801), .FEN(FEN[3551]), .op(N5801_t1) );
fim FAN_N5798_0 ( .fault(fault), .net(N5798), .FEN(FEN[3552]), .op(N5798_t0) );
fim FAN_N5798_1 ( .fault(fault), .net(N5798), .FEN(FEN[3553]), .op(N5798_t1) );
fim FAN_N5804_0 ( .fault(fault), .net(N5804), .FEN(FEN[3554]), .op(N5804_t0) );
fim FAN_N5804_1 ( .fault(fault), .net(N5804), .FEN(FEN[3555]), .op(N5804_t1) );
fim FAN_N5804_2 ( .fault(fault), .net(N5804), .FEN(FEN[3556]), .op(N5804_t2) );
fim FAN_N5810_0 ( .fault(fault), .net(N5810), .FEN(FEN[3557]), .op(N5810_t0) );
fim FAN_N5810_1 ( .fault(fault), .net(N5810), .FEN(FEN[3558]), .op(N5810_t1) );
fim FAN_N924_0 ( .fault(fault), .net(N924), .FEN(FEN[3559]), .op(N924_t0) );
fim FAN_N924_1 ( .fault(fault), .net(N924), .FEN(FEN[3560]), .op(N924_t1) );
fim FAN_N5813_0 ( .fault(fault), .net(N5813), .FEN(FEN[3561]), .op(N5813_t0) );
fim FAN_N5813_1 ( .fault(fault), .net(N5813), .FEN(FEN[3562]), .op(N5813_t1) );
fim FAN_N5813_2 ( .fault(fault), .net(N5813), .FEN(FEN[3563]), .op(N5813_t2) );
fim FAN_N5822_0 ( .fault(fault), .net(N5822), .FEN(FEN[3564]), .op(N5822_t0) );
fim FAN_N5822_1 ( .fault(fault), .net(N5822), .FEN(FEN[3565]), .op(N5822_t1) );
fim FAN_N5819_0 ( .fault(fault), .net(N5819), .FEN(FEN[3566]), .op(N5819_t0) );
fim FAN_N5819_1 ( .fault(fault), .net(N5819), .FEN(FEN[3567]), .op(N5819_t1) );
fim FAN_N5825_0 ( .fault(fault), .net(N5825), .FEN(FEN[3568]), .op(N5825_t0) );
fim FAN_N5825_1 ( .fault(fault), .net(N5825), .FEN(FEN[3569]), .op(N5825_t1) );
fim FAN_N5825_2 ( .fault(fault), .net(N5825), .FEN(FEN[3570]), .op(N5825_t2) );
fim FAN_N5834_0 ( .fault(fault), .net(N5834), .FEN(FEN[3571]), .op(N5834_t0) );
fim FAN_N5834_1 ( .fault(fault), .net(N5834), .FEN(FEN[3572]), .op(N5834_t1) );
fim FAN_N585_0 ( .fault(fault), .net(N585), .FEN(FEN[3573]), .op(N585_t0) );
fim FAN_N585_1 ( .fault(fault), .net(N585), .FEN(FEN[3574]), .op(N585_t1) );
fim FAN_N5837_0 ( .fault(fault), .net(N5837), .FEN(FEN[3575]), .op(N5837_t0) );
fim FAN_N5837_1 ( .fault(fault), .net(N5837), .FEN(FEN[3576]), .op(N5837_t1) );
fim FAN_N633_0 ( .fault(fault), .net(N633), .FEN(FEN[3577]), .op(N633_t0) );
fim FAN_N633_1 ( .fault(fault), .net(N633), .FEN(FEN[3578]), .op(N633_t1) );
fim FAN_N5840_0 ( .fault(fault), .net(N5840), .FEN(FEN[3579]), .op(N5840_t0) );
fim FAN_N5840_1 ( .fault(fault), .net(N5840), .FEN(FEN[3580]), .op(N5840_t1) );
fim FAN_N5840_2 ( .fault(fault), .net(N5840), .FEN(FEN[3581]), .op(N5840_t2) );
fim FAN_N5849_0 ( .fault(fault), .net(N5849), .FEN(FEN[3582]), .op(N5849_t0) );
fim FAN_N5849_1 ( .fault(fault), .net(N5849), .FEN(FEN[3583]), .op(N5849_t1) );
fim FAN_N5846_0 ( .fault(fault), .net(N5846), .FEN(FEN[3584]), .op(N5846_t0) );
fim FAN_N5846_1 ( .fault(fault), .net(N5846), .FEN(FEN[3585]), .op(N5846_t1) );
fim FAN_N5852_0 ( .fault(fault), .net(N5852), .FEN(FEN[3586]), .op(N5852_t0) );
fim FAN_N5852_1 ( .fault(fault), .net(N5852), .FEN(FEN[3587]), .op(N5852_t1) );
fim FAN_N5852_2 ( .fault(fault), .net(N5852), .FEN(FEN[3588]), .op(N5852_t2) );
fim FAN_N5858_0 ( .fault(fault), .net(N5858), .FEN(FEN[3589]), .op(N5858_t0) );
fim FAN_N5858_1 ( .fault(fault), .net(N5858), .FEN(FEN[3590]), .op(N5858_t1) );
fim FAN_N876_0 ( .fault(fault), .net(N876), .FEN(FEN[3591]), .op(N876_t0) );
fim FAN_N876_1 ( .fault(fault), .net(N876), .FEN(FEN[3592]), .op(N876_t1) );
fim FAN_N5861_0 ( .fault(fault), .net(N5861), .FEN(FEN[3593]), .op(N5861_t0) );
fim FAN_N5861_1 ( .fault(fault), .net(N5861), .FEN(FEN[3594]), .op(N5861_t1) );
fim FAN_N5861_2 ( .fault(fault), .net(N5861), .FEN(FEN[3595]), .op(N5861_t2) );
fim FAN_N5870_0 ( .fault(fault), .net(N5870), .FEN(FEN[3596]), .op(N5870_t0) );
fim FAN_N5870_1 ( .fault(fault), .net(N5870), .FEN(FEN[3597]), .op(N5870_t1) );
fim FAN_N5867_0 ( .fault(fault), .net(N5867), .FEN(FEN[3598]), .op(N5867_t0) );
fim FAN_N5867_1 ( .fault(fault), .net(N5867), .FEN(FEN[3599]), .op(N5867_t1) );
fim FAN_N5873_0 ( .fault(fault), .net(N5873), .FEN(FEN[3600]), .op(N5873_t0) );
fim FAN_N5873_1 ( .fault(fault), .net(N5873), .FEN(FEN[3601]), .op(N5873_t1) );
fim FAN_N5873_2 ( .fault(fault), .net(N5873), .FEN(FEN[3602]), .op(N5873_t2) );
fim FAN_N5882_0 ( .fault(fault), .net(N5882), .FEN(FEN[3603]), .op(N5882_t0) );
fim FAN_N5882_1 ( .fault(fault), .net(N5882), .FEN(FEN[3604]), .op(N5882_t1) );
fim FAN_N5882_2 ( .fault(fault), .net(N5882), .FEN(FEN[3605]), .op(N5882_t2) );
fim FAN_N5886_0 ( .fault(fault), .net(N5886), .FEN(FEN[3606]), .op(N5886_t0) );
fim FAN_N5886_1 ( .fault(fault), .net(N5886), .FEN(FEN[3607]), .op(N5886_t1) );
fim FAN_N5886_2 ( .fault(fault), .net(N5886), .FEN(FEN[3608]), .op(N5886_t2) );
fim FAN_N5895_0 ( .fault(fault), .net(N5895), .FEN(FEN[3609]), .op(N5895_t0) );
fim FAN_N5895_1 ( .fault(fault), .net(N5895), .FEN(FEN[3610]), .op(N5895_t1) );
fim FAN_N5892_0 ( .fault(fault), .net(N5892), .FEN(FEN[3611]), .op(N5892_t0) );
fim FAN_N5892_1 ( .fault(fault), .net(N5892), .FEN(FEN[3612]), .op(N5892_t1) );
fim FAN_N5898_0 ( .fault(fault), .net(N5898), .FEN(FEN[3613]), .op(N5898_t0) );
fim FAN_N5898_1 ( .fault(fault), .net(N5898), .FEN(FEN[3614]), .op(N5898_t1) );
fim FAN_N5898_2 ( .fault(fault), .net(N5898), .FEN(FEN[3615]), .op(N5898_t2) );
fim FAN_N5904_0 ( .fault(fault), .net(N5904), .FEN(FEN[3616]), .op(N5904_t0) );
fim FAN_N5904_1 ( .fault(fault), .net(N5904), .FEN(FEN[3617]), .op(N5904_t1) );
fim FAN_N828_0 ( .fault(fault), .net(N828), .FEN(FEN[3618]), .op(N828_t0) );
fim FAN_N828_1 ( .fault(fault), .net(N828), .FEN(FEN[3619]), .op(N828_t1) );
fim FAN_N5907_0 ( .fault(fault), .net(N5907), .FEN(FEN[3620]), .op(N5907_t0) );
fim FAN_N5907_1 ( .fault(fault), .net(N5907), .FEN(FEN[3621]), .op(N5907_t1) );
fim FAN_N5907_2 ( .fault(fault), .net(N5907), .FEN(FEN[3622]), .op(N5907_t2) );
fim FAN_N5916_0 ( .fault(fault), .net(N5916), .FEN(FEN[3623]), .op(N5916_t0) );
fim FAN_N5916_1 ( .fault(fault), .net(N5916), .FEN(FEN[3624]), .op(N5916_t1) );
fim FAN_N5913_0 ( .fault(fault), .net(N5913), .FEN(FEN[3625]), .op(N5913_t0) );
fim FAN_N5913_1 ( .fault(fault), .net(N5913), .FEN(FEN[3626]), .op(N5913_t1) );
fim FAN_N5919_0 ( .fault(fault), .net(N5919), .FEN(FEN[3627]), .op(N5919_t0) );
fim FAN_N5919_1 ( .fault(fault), .net(N5919), .FEN(FEN[3628]), .op(N5919_t1) );
fim FAN_N5919_2 ( .fault(fault), .net(N5919), .FEN(FEN[3629]), .op(N5919_t2) );
fim FAN_N5938_0 ( .fault(fault), .net(N5938), .FEN(FEN[3630]), .op(N5938_t0) );
fim FAN_N5938_1 ( .fault(fault), .net(N5938), .FEN(FEN[3631]), .op(N5938_t1) );
fim FAN_N5935_0 ( .fault(fault), .net(N5935), .FEN(FEN[3632]), .op(N5935_t0) );
fim FAN_N5935_1 ( .fault(fault), .net(N5935), .FEN(FEN[3633]), .op(N5935_t1) );
fim FAN_N5941_0 ( .fault(fault), .net(N5941), .FEN(FEN[3634]), .op(N5941_t0) );
fim FAN_N5941_1 ( .fault(fault), .net(N5941), .FEN(FEN[3635]), .op(N5941_t1) );
fim FAN_N5941_2 ( .fault(fault), .net(N5941), .FEN(FEN[3636]), .op(N5941_t2) );
fim FAN_N5947_0 ( .fault(fault), .net(N5947), .FEN(FEN[3637]), .op(N5947_t0) );
fim FAN_N5947_1 ( .fault(fault), .net(N5947), .FEN(FEN[3638]), .op(N5947_t1) );
fim FAN_N780_0 ( .fault(fault), .net(N780), .FEN(FEN[3639]), .op(N780_t0) );
fim FAN_N780_1 ( .fault(fault), .net(N780), .FEN(FEN[3640]), .op(N780_t1) );
fim FAN_N5950_0 ( .fault(fault), .net(N5950), .FEN(FEN[3641]), .op(N5950_t0) );
fim FAN_N5950_1 ( .fault(fault), .net(N5950), .FEN(FEN[3642]), .op(N5950_t1) );
fim FAN_N5950_2 ( .fault(fault), .net(N5950), .FEN(FEN[3643]), .op(N5950_t2) );
fim FAN_N5959_0 ( .fault(fault), .net(N5959), .FEN(FEN[3644]), .op(N5959_t0) );
fim FAN_N5959_1 ( .fault(fault), .net(N5959), .FEN(FEN[3645]), .op(N5959_t1) );
fim FAN_N5956_0 ( .fault(fault), .net(N5956), .FEN(FEN[3646]), .op(N5956_t0) );
fim FAN_N5956_1 ( .fault(fault), .net(N5956), .FEN(FEN[3647]), .op(N5956_t1) );
fim FAN_N5962_0 ( .fault(fault), .net(N5962), .FEN(FEN[3648]), .op(N5962_t0) );
fim FAN_N5962_1 ( .fault(fault), .net(N5962), .FEN(FEN[3649]), .op(N5962_t1) );
fim FAN_N5962_2 ( .fault(fault), .net(N5962), .FEN(FEN[3650]), .op(N5962_t2) );
fim FAN_N5972_0 ( .fault(fault), .net(N5972), .FEN(FEN[3651]), .op(N5972_t0) );
fim FAN_N5972_1 ( .fault(fault), .net(N5972), .FEN(FEN[3652]), .op(N5972_t1) );
fim FAN_N5930_0 ( .fault(fault), .net(N5930), .FEN(FEN[3653]), .op(N5930_t0) );
fim FAN_N5930_1 ( .fault(fault), .net(N5930), .FEN(FEN[3654]), .op(N5930_t1) );
fim FAN_N5975_0 ( .fault(fault), .net(N5975), .FEN(FEN[3655]), .op(N5975_t0) );
fim FAN_N5975_1 ( .fault(fault), .net(N5975), .FEN(FEN[3656]), .op(N5975_t1) );
fim FAN_N5975_2 ( .fault(fault), .net(N5975), .FEN(FEN[3657]), .op(N5975_t2) );
fim FAN_N5981_0 ( .fault(fault), .net(N5981), .FEN(FEN[3658]), .op(N5981_t0) );
fim FAN_N5981_1 ( .fault(fault), .net(N5981), .FEN(FEN[3659]), .op(N5981_t1) );
fim FAN_N732_0 ( .fault(fault), .net(N732), .FEN(FEN[3660]), .op(N732_t0) );
fim FAN_N732_1 ( .fault(fault), .net(N732), .FEN(FEN[3661]), .op(N732_t1) );
fim FAN_N5984_0 ( .fault(fault), .net(N5984), .FEN(FEN[3662]), .op(N5984_t0) );
fim FAN_N5984_1 ( .fault(fault), .net(N5984), .FEN(FEN[3663]), .op(N5984_t1) );
fim FAN_N5984_2 ( .fault(fault), .net(N5984), .FEN(FEN[3664]), .op(N5984_t2) );
fim FAN_N5993_0 ( .fault(fault), .net(N5993), .FEN(FEN[3665]), .op(N5993_t0) );
fim FAN_N5993_1 ( .fault(fault), .net(N5993), .FEN(FEN[3666]), .op(N5993_t1) );
fim FAN_N5990_0 ( .fault(fault), .net(N5990), .FEN(FEN[3667]), .op(N5990_t0) );
fim FAN_N5990_1 ( .fault(fault), .net(N5990), .FEN(FEN[3668]), .op(N5990_t1) );
fim FAN_N5996_0 ( .fault(fault), .net(N5996), .FEN(FEN[3669]), .op(N5996_t0) );
fim FAN_N5996_1 ( .fault(fault), .net(N5996), .FEN(FEN[3670]), .op(N5996_t1) );
fim FAN_N5996_2 ( .fault(fault), .net(N5996), .FEN(FEN[3671]), .op(N5996_t2) );
fim FAN_N6005_0 ( .fault(fault), .net(N6005), .FEN(FEN[3672]), .op(N6005_t0) );
fim FAN_N6005_1 ( .fault(fault), .net(N6005), .FEN(FEN[3673]), .op(N6005_t1) );
fim FAN_N6005_2 ( .fault(fault), .net(N6005), .FEN(FEN[3674]), .op(N6005_t2) );
fim FAN_N6011_0 ( .fault(fault), .net(N6011), .FEN(FEN[3675]), .op(N6011_t0) );
fim FAN_N6011_1 ( .fault(fault), .net(N6011), .FEN(FEN[3676]), .op(N6011_t1) );
fim FAN_N684_0 ( .fault(fault), .net(N684), .FEN(FEN[3677]), .op(N684_t0) );
fim FAN_N684_1 ( .fault(fault), .net(N684), .FEN(FEN[3678]), .op(N684_t1) );
fim FAN_N6014_0 ( .fault(fault), .net(N6014), .FEN(FEN[3679]), .op(N6014_t0) );
fim FAN_N6014_1 ( .fault(fault), .net(N6014), .FEN(FEN[3680]), .op(N6014_t1) );
fim FAN_N6014_2 ( .fault(fault), .net(N6014), .FEN(FEN[3681]), .op(N6014_t2) );
fim FAN_N6023_0 ( .fault(fault), .net(N6023), .FEN(FEN[3682]), .op(N6023_t0) );
fim FAN_N6023_1 ( .fault(fault), .net(N6023), .FEN(FEN[3683]), .op(N6023_t1) );
fim FAN_N6020_0 ( .fault(fault), .net(N6020), .FEN(FEN[3684]), .op(N6020_t0) );
fim FAN_N6020_1 ( .fault(fault), .net(N6020), .FEN(FEN[3685]), .op(N6020_t1) );
fim FAN_N6026_0 ( .fault(fault), .net(N6026), .FEN(FEN[3686]), .op(N6026_t0) );
fim FAN_N6026_1 ( .fault(fault), .net(N6026), .FEN(FEN[3687]), .op(N6026_t1) );
fim FAN_N6026_2 ( .fault(fault), .net(N6026), .FEN(FEN[3688]), .op(N6026_t2) );
fim FAN_N6037_0 ( .fault(fault), .net(N6037), .FEN(FEN[3689]), .op(N6037_t0) );
fim FAN_N6037_1 ( .fault(fault), .net(N6037), .FEN(FEN[3690]), .op(N6037_t1) );
fim FAN_N636_0 ( .fault(fault), .net(N636), .FEN(FEN[3691]), .op(N636_t0) );
fim FAN_N636_1 ( .fault(fault), .net(N636), .FEN(FEN[3692]), .op(N636_t1) );
fim FAN_N6040_0 ( .fault(fault), .net(N6040), .FEN(FEN[3693]), .op(N6040_t0) );
fim FAN_N6040_1 ( .fault(fault), .net(N6040), .FEN(FEN[3694]), .op(N6040_t1) );
fim FAN_N6040_2 ( .fault(fault), .net(N6040), .FEN(FEN[3695]), .op(N6040_t2) );
fim FAN_N6049_0 ( .fault(fault), .net(N6049), .FEN(FEN[3696]), .op(N6049_t0) );
fim FAN_N6049_1 ( .fault(fault), .net(N6049), .FEN(FEN[3697]), .op(N6049_t1) );
fim FAN_N6046_0 ( .fault(fault), .net(N6046), .FEN(FEN[3698]), .op(N6046_t0) );
fim FAN_N6046_1 ( .fault(fault), .net(N6046), .FEN(FEN[3699]), .op(N6046_t1) );
fim FAN_N6052_0 ( .fault(fault), .net(N6052), .FEN(FEN[3700]), .op(N6052_t0) );
fim FAN_N6052_1 ( .fault(fault), .net(N6052), .FEN(FEN[3701]), .op(N6052_t1) );
fim FAN_N6052_2 ( .fault(fault), .net(N6052), .FEN(FEN[3702]), .op(N6052_t2) );
fim FAN_N6061_0 ( .fault(fault), .net(N6061), .FEN(FEN[3703]), .op(N6061_t0) );
fim FAN_N6061_1 ( .fault(fault), .net(N6061), .FEN(FEN[3704]), .op(N6061_t1) );
fim FAN_N588_0 ( .fault(fault), .net(N588), .FEN(FEN[3705]), .op(N588_t0) );
fim FAN_N588_1 ( .fault(fault), .net(N588), .FEN(FEN[3706]), .op(N588_t1) );
fim FAN_N6064_0 ( .fault(fault), .net(N6064), .FEN(FEN[3707]), .op(N6064_t0) );
fim FAN_N6064_1 ( .fault(fault), .net(N6064), .FEN(FEN[3708]), .op(N6064_t1) );
fim FAN_N6064_2 ( .fault(fault), .net(N6064), .FEN(FEN[3709]), .op(N6064_t2) );
fim FAN_N6073_0 ( .fault(fault), .net(N6073), .FEN(FEN[3710]), .op(N6073_t0) );
fim FAN_N6073_1 ( .fault(fault), .net(N6073), .FEN(FEN[3711]), .op(N6073_t1) );
fim FAN_N6070_0 ( .fault(fault), .net(N6070), .FEN(FEN[3712]), .op(N6070_t0) );
fim FAN_N6070_1 ( .fault(fault), .net(N6070), .FEN(FEN[3713]), .op(N6070_t1) );
fim FAN_N6076_0 ( .fault(fault), .net(N6076), .FEN(FEN[3714]), .op(N6076_t0) );
fim FAN_N6076_1 ( .fault(fault), .net(N6076), .FEN(FEN[3715]), .op(N6076_t1) );
fim FAN_N6076_2 ( .fault(fault), .net(N6076), .FEN(FEN[3716]), .op(N6076_t2) );
fim FAN_N6085_0 ( .fault(fault), .net(N6085), .FEN(FEN[3717]), .op(N6085_t0) );
fim FAN_N6085_1 ( .fault(fault), .net(N6085), .FEN(FEN[3718]), .op(N6085_t1) );
fim FAN_N6085_2 ( .fault(fault), .net(N6085), .FEN(FEN[3719]), .op(N6085_t2) );
fim FAN_N6094_0 ( .fault(fault), .net(N6094), .FEN(FEN[3720]), .op(N6094_t0) );
fim FAN_N6094_1 ( .fault(fault), .net(N6094), .FEN(FEN[3721]), .op(N6094_t1) );
fim FAN_N6091_0 ( .fault(fault), .net(N6091), .FEN(FEN[3722]), .op(N6091_t0) );
fim FAN_N6091_1 ( .fault(fault), .net(N6091), .FEN(FEN[3723]), .op(N6091_t1) );
fim FAN_N6097_0 ( .fault(fault), .net(N6097), .FEN(FEN[3724]), .op(N6097_t0) );
fim FAN_N6097_1 ( .fault(fault), .net(N6097), .FEN(FEN[3725]), .op(N6097_t1) );
fim FAN_N6097_2 ( .fault(fault), .net(N6097), .FEN(FEN[3726]), .op(N6097_t2) );
fim FAN_N6111_0 ( .fault(fault), .net(N6111), .FEN(FEN[3727]), .op(N6111_t0) );
fim FAN_N6111_1 ( .fault(fault), .net(N6111), .FEN(FEN[3728]), .op(N6111_t1) );
fim FAN_N6108_0 ( .fault(fault), .net(N6108), .FEN(FEN[3729]), .op(N6108_t0) );
fim FAN_N6108_1 ( .fault(fault), .net(N6108), .FEN(FEN[3730]), .op(N6108_t1) );
fim FAN_N6114_0 ( .fault(fault), .net(N6114), .FEN(FEN[3731]), .op(N6114_t0) );
fim FAN_N6114_1 ( .fault(fault), .net(N6114), .FEN(FEN[3732]), .op(N6114_t1) );
fim FAN_N6114_2 ( .fault(fault), .net(N6114), .FEN(FEN[3733]), .op(N6114_t2) );
fim FAN_N6124_0 ( .fault(fault), .net(N6124), .FEN(FEN[3734]), .op(N6124_t0) );
fim FAN_N6124_1 ( .fault(fault), .net(N6124), .FEN(FEN[3735]), .op(N6124_t1) );
fim FAN_N6124_2 ( .fault(fault), .net(N6124), .FEN(FEN[3736]), .op(N6124_t2) );
fim FAN_N6138_0 ( .fault(fault), .net(N6138), .FEN(FEN[3737]), .op(N6138_t0) );
fim FAN_N6138_1 ( .fault(fault), .net(N6138), .FEN(FEN[3738]), .op(N6138_t1) );
fim FAN_N6141_0 ( .fault(fault), .net(N6141), .FEN(FEN[3739]), .op(N6141_t0) );
fim FAN_N6141_1 ( .fault(fault), .net(N6141), .FEN(FEN[3740]), .op(N6141_t1) );
fim FAN_N6141_2 ( .fault(fault), .net(N6141), .FEN(FEN[3741]), .op(N6141_t2) );
fim FAN_N6135_0 ( .fault(fault), .net(N6135), .FEN(FEN[3742]), .op(N6135_t0) );
fim FAN_N6135_1 ( .fault(fault), .net(N6135), .FEN(FEN[3743]), .op(N6135_t1) );
fim FAN_N6147_0 ( .fault(fault), .net(N6147), .FEN(FEN[3744]), .op(N6147_t0) );
fim FAN_N6147_1 ( .fault(fault), .net(N6147), .FEN(FEN[3745]), .op(N6147_t1) );
fim FAN_N6151_0 ( .fault(fault), .net(N6151), .FEN(FEN[3746]), .op(N6151_t0) );
fim FAN_N6151_1 ( .fault(fault), .net(N6151), .FEN(FEN[3747]), .op(N6151_t1) );
fim FAN_N6151_2 ( .fault(fault), .net(N6151), .FEN(FEN[3748]), .op(N6151_t2) );
fim FAN_N6130_0 ( .fault(fault), .net(N6130), .FEN(FEN[3749]), .op(N6130_t0) );
fim FAN_N6130_1 ( .fault(fault), .net(N6130), .FEN(FEN[3750]), .op(N6130_t1) );
fim FAN_N6157_0 ( .fault(fault), .net(N6157), .FEN(FEN[3751]), .op(N6157_t0) );
fim FAN_N6157_1 ( .fault(fault), .net(N6157), .FEN(FEN[3752]), .op(N6157_t1) );
fim FAN_N6161_0 ( .fault(fault), .net(N6161), .FEN(FEN[3753]), .op(N6161_t0) );
fim FAN_N6161_1 ( .fault(fault), .net(N6161), .FEN(FEN[3754]), .op(N6161_t1) );
fim FAN_N6161_2 ( .fault(fault), .net(N6161), .FEN(FEN[3755]), .op(N6161_t2) );
fim FAN_N6120_0 ( .fault(fault), .net(N6120), .FEN(FEN[3756]), .op(N6120_t0) );
fim FAN_N6120_1 ( .fault(fault), .net(N6120), .FEN(FEN[3757]), .op(N6120_t1) );
fim FAN_N6167_0 ( .fault(fault), .net(N6167), .FEN(FEN[3758]), .op(N6167_t0) );
fim FAN_N6167_1 ( .fault(fault), .net(N6167), .FEN(FEN[3759]), .op(N6167_t1) );
fim FAN_N6171_0 ( .fault(fault), .net(N6171), .FEN(FEN[3760]), .op(N6171_t0) );
fim FAN_N6171_1 ( .fault(fault), .net(N6171), .FEN(FEN[3761]), .op(N6171_t1) );
fim FAN_N6171_2 ( .fault(fault), .net(N6171), .FEN(FEN[3762]), .op(N6171_t2) );
fim FAN_N6103_0 ( .fault(fault), .net(N6103), .FEN(FEN[3763]), .op(N6103_t0) );
fim FAN_N6103_1 ( .fault(fault), .net(N6103), .FEN(FEN[3764]), .op(N6103_t1) );
fim FAN_N6177_0 ( .fault(fault), .net(N6177), .FEN(FEN[3765]), .op(N6177_t0) );
fim FAN_N6177_1 ( .fault(fault), .net(N6177), .FEN(FEN[3766]), .op(N6177_t1) );
fim FAN_N6181_0 ( .fault(fault), .net(N6181), .FEN(FEN[3767]), .op(N6181_t0) );
fim FAN_N6181_1 ( .fault(fault), .net(N6181), .FEN(FEN[3768]), .op(N6181_t1) );
fim FAN_N6181_2 ( .fault(fault), .net(N6181), .FEN(FEN[3769]), .op(N6181_t2) );
fim FAN_N6082_0 ( .fault(fault), .net(N6082), .FEN(FEN[3770]), .op(N6082_t0) );
fim FAN_N6082_1 ( .fault(fault), .net(N6082), .FEN(FEN[3771]), .op(N6082_t1) );
fim FAN_N6187_0 ( .fault(fault), .net(N6187), .FEN(FEN[3772]), .op(N6187_t0) );
fim FAN_N6187_1 ( .fault(fault), .net(N6187), .FEN(FEN[3773]), .op(N6187_t1) );
fim FAN_N6191_0 ( .fault(fault), .net(N6191), .FEN(FEN[3774]), .op(N6191_t0) );
fim FAN_N6191_1 ( .fault(fault), .net(N6191), .FEN(FEN[3775]), .op(N6191_t1) );
fim FAN_N6191_2 ( .fault(fault), .net(N6191), .FEN(FEN[3776]), .op(N6191_t2) );
fim FAN_N6058_0 ( .fault(fault), .net(N6058), .FEN(FEN[3777]), .op(N6058_t0) );
fim FAN_N6058_1 ( .fault(fault), .net(N6058), .FEN(FEN[3778]), .op(N6058_t1) );
fim FAN_N6197_0 ( .fault(fault), .net(N6197), .FEN(FEN[3779]), .op(N6197_t0) );
fim FAN_N6197_1 ( .fault(fault), .net(N6197), .FEN(FEN[3780]), .op(N6197_t1) );
fim FAN_N6201_0 ( .fault(fault), .net(N6201), .FEN(FEN[3781]), .op(N6201_t0) );
fim FAN_N6201_1 ( .fault(fault), .net(N6201), .FEN(FEN[3782]), .op(N6201_t1) );
fim FAN_N6201_2 ( .fault(fault), .net(N6201), .FEN(FEN[3783]), .op(N6201_t2) );
fim FAN_N6032_0 ( .fault(fault), .net(N6032), .FEN(FEN[3784]), .op(N6032_t0) );
fim FAN_N6032_1 ( .fault(fault), .net(N6032), .FEN(FEN[3785]), .op(N6032_t1) );
fim FAN_N6207_0 ( .fault(fault), .net(N6207), .FEN(FEN[3786]), .op(N6207_t0) );
fim FAN_N6207_1 ( .fault(fault), .net(N6207), .FEN(FEN[3787]), .op(N6207_t1) );
fim FAN_N6211_0 ( .fault(fault), .net(N6211), .FEN(FEN[3788]), .op(N6211_t0) );
fim FAN_N6211_1 ( .fault(fault), .net(N6211), .FEN(FEN[3789]), .op(N6211_t1) );
fim FAN_N6211_2 ( .fault(fault), .net(N6211), .FEN(FEN[3790]), .op(N6211_t2) );
fim FAN_N6002_0 ( .fault(fault), .net(N6002), .FEN(FEN[3791]), .op(N6002_t0) );
fim FAN_N6002_1 ( .fault(fault), .net(N6002), .FEN(FEN[3792]), .op(N6002_t1) );
fim FAN_N6217_0 ( .fault(fault), .net(N6217), .FEN(FEN[3793]), .op(N6217_t0) );
fim FAN_N6217_1 ( .fault(fault), .net(N6217), .FEN(FEN[3794]), .op(N6217_t1) );
fim FAN_N6221_0 ( .fault(fault), .net(N6221), .FEN(FEN[3795]), .op(N6221_t0) );
fim FAN_N6221_1 ( .fault(fault), .net(N6221), .FEN(FEN[3796]), .op(N6221_t1) );
fim FAN_N6221_2 ( .fault(fault), .net(N6221), .FEN(FEN[3797]), .op(N6221_t2) );
fim FAN_N5968_0 ( .fault(fault), .net(N5968), .FEN(FEN[3798]), .op(N5968_t0) );
fim FAN_N5968_1 ( .fault(fault), .net(N5968), .FEN(FEN[3799]), .op(N5968_t1) );
fim FAN_N6227_0 ( .fault(fault), .net(N6227), .FEN(FEN[3800]), .op(N6227_t0) );
fim FAN_N6227_1 ( .fault(fault), .net(N6227), .FEN(FEN[3801]), .op(N6227_t1) );
fim FAN_N6231_0 ( .fault(fault), .net(N6231), .FEN(FEN[3802]), .op(N6231_t0) );
fim FAN_N6231_1 ( .fault(fault), .net(N6231), .FEN(FEN[3803]), .op(N6231_t1) );
fim FAN_N6231_2 ( .fault(fault), .net(N6231), .FEN(FEN[3804]), .op(N6231_t2) );
fim FAN_N5925_0 ( .fault(fault), .net(N5925), .FEN(FEN[3805]), .op(N5925_t0) );
fim FAN_N5925_1 ( .fault(fault), .net(N5925), .FEN(FEN[3806]), .op(N5925_t1) );
fim FAN_N6237_0 ( .fault(fault), .net(N6237), .FEN(FEN[3807]), .op(N6237_t0) );
fim FAN_N6237_1 ( .fault(fault), .net(N6237), .FEN(FEN[3808]), .op(N6237_t1) );
fim FAN_N6241_0 ( .fault(fault), .net(N6241), .FEN(FEN[3809]), .op(N6241_t0) );
fim FAN_N6241_1 ( .fault(fault), .net(N6241), .FEN(FEN[3810]), .op(N6241_t1) );
fim FAN_N6241_2 ( .fault(fault), .net(N6241), .FEN(FEN[3811]), .op(N6241_t2) );
fim FAN_N5879_0 ( .fault(fault), .net(N5879), .FEN(FEN[3812]), .op(N5879_t0) );
fim FAN_N5879_1 ( .fault(fault), .net(N5879), .FEN(FEN[3813]), .op(N5879_t1) );
fim FAN_N6247_0 ( .fault(fault), .net(N6247), .FEN(FEN[3814]), .op(N6247_t0) );
fim FAN_N6247_1 ( .fault(fault), .net(N6247), .FEN(FEN[3815]), .op(N6247_t1) );
fim FAN_N6251_0 ( .fault(fault), .net(N6251), .FEN(FEN[3816]), .op(N6251_t0) );
fim FAN_N6251_1 ( .fault(fault), .net(N6251), .FEN(FEN[3817]), .op(N6251_t1) );
fim FAN_N6251_2 ( .fault(fault), .net(N6251), .FEN(FEN[3818]), .op(N6251_t2) );
fim FAN_N5831_0 ( .fault(fault), .net(N5831), .FEN(FEN[3819]), .op(N5831_t0) );
fim FAN_N5831_1 ( .fault(fault), .net(N5831), .FEN(FEN[3820]), .op(N5831_t1) );
fim FAN_N6257_0 ( .fault(fault), .net(N6257), .FEN(FEN[3821]), .op(N6257_t0) );
fim FAN_N6257_1 ( .fault(fault), .net(N6257), .FEN(FEN[3822]), .op(N6257_t1) );
fim FAN_N6261_0 ( .fault(fault), .net(N6261), .FEN(FEN[3823]), .op(N6261_t0) );
fim FAN_N6261_1 ( .fault(fault), .net(N6261), .FEN(FEN[3824]), .op(N6261_t1) );
fim FAN_N6261_2 ( .fault(fault), .net(N6261), .FEN(FEN[3825]), .op(N6261_t2) );
fim FAN_N5782_0 ( .fault(fault), .net(N5782), .FEN(FEN[3826]), .op(N5782_t0) );
fim FAN_N5782_1 ( .fault(fault), .net(N5782), .FEN(FEN[3827]), .op(N5782_t1) );
fim FAN_N6267_0 ( .fault(fault), .net(N6267), .FEN(FEN[3828]), .op(N6267_t0) );
fim FAN_N6267_1 ( .fault(fault), .net(N6267), .FEN(FEN[3829]), .op(N6267_t1) );
fim FAN_N6271_0 ( .fault(fault), .net(N6271), .FEN(FEN[3830]), .op(N6271_t0) );
fim FAN_N6271_1 ( .fault(fault), .net(N6271), .FEN(FEN[3831]), .op(N6271_t1) );
fim FAN_N6271_2 ( .fault(fault), .net(N6271), .FEN(FEN[3832]), .op(N6271_t2) );
fim FAN_N5727_0 ( .fault(fault), .net(N5727), .FEN(FEN[3833]), .op(N5727_t0) );
fim FAN_N5727_1 ( .fault(fault), .net(N5727), .FEN(FEN[3834]), .op(N5727_t1) );
fim FAN_N6277_0 ( .fault(fault), .net(N6277), .FEN(FEN[3835]), .op(N6277_t0) );
fim FAN_N6277_1 ( .fault(fault), .net(N6277), .FEN(FEN[3836]), .op(N6277_t1) );
fim FAN_N6281_0 ( .fault(fault), .net(N6281), .FEN(FEN[3837]), .op(N6281_t0) );
fim FAN_N6281_1 ( .fault(fault), .net(N6281), .FEN(FEN[3838]), .op(N6281_t1) );
fim FAN_N6281_2 ( .fault(fault), .net(N6281), .FEN(FEN[3839]), .op(N6281_t2) );
initial begin
    FEN <= {3839'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {3839'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,3839'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,3839'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN <= {FEN[3838:0], FEN[3839]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
// EndFaultModel

//Anchor
and AND2_1 (N545, N1_t0, N273_t0);
and AND2_2 (N546, N1_t1, N290_t0);
and AND2_3 (N549, N1_t2, N307_t0);
and AND2_4 (N552, N1_t3, N324_t0);
and AND2_5 (N555, N1_t4, N341_t0);
and AND2_6 (N558, N1_t5, N358_t0);
and AND2_7 (N561, N1_t6, N375_t0);
and AND2_8 (N564, N1_t7, N392_t0);
and AND2_9 (N567, N1_t8, N409_t0);
and AND2_10 (N570, N1_t9, N426_t0);
and AND2_11 (N573, N1_t10, N443_t0);
and AND2_12 (N576, N1_t11, N460_t0);
and AND2_13 (N579, N1_t12, N477_t0);
and AND2_14 (N582, N1_t13, N494_t0);
and AND2_15 (N585, N1_t14, N511_t0);
and AND2_16 (N588, N1_t15, N528_t0);
and AND2_17 (N591, N18_t0, N273_t1);
and AND2_18 (N594, N18_t1, N290_t1);
and AND2_19 (N597, N18_t2, N307_t1);
and AND2_20 (N600, N18_t3, N324_t1);
and AND2_21 (N603, N18_t4, N341_t1);
and AND2_22 (N606, N18_t5, N358_t1);
and AND2_23 (N609, N18_t6, N375_t1);
and AND2_24 (N612, N18_t7, N392_t1);
and AND2_25 (N615, N18_t8, N409_t1);
and AND2_26 (N618, N18_t9, N426_t1);
and AND2_27 (N621, N18_t10, N443_t1);
and AND2_28 (N624, N18_t11, N460_t1);
and AND2_29 (N627, N18_t12, N477_t1);
and AND2_30 (N630, N18_t13, N494_t1);
and AND2_31 (N633, N18_t14, N511_t1);
and AND2_32 (N636, N18_t15, N528_t1);
and AND2_33 (N639, N35_t0, N273_t2);
and AND2_34 (N642, N35_t1, N290_t2);
and AND2_35 (N645, N35_t2, N307_t2);
and AND2_36 (N648, N35_t3, N324_t2);
and AND2_37 (N651, N35_t4, N341_t2);
and AND2_38 (N654, N35_t5, N358_t2);
and AND2_39 (N657, N35_t6, N375_t2);
and AND2_40 (N660, N35_t7, N392_t2);
and AND2_41 (N663, N35_t8, N409_t2);
and AND2_42 (N666, N35_t9, N426_t2);
and AND2_43 (N669, N35_t10, N443_t2);
and AND2_44 (N672, N35_t11, N460_t2);
and AND2_45 (N675, N35_t12, N477_t2);
and AND2_46 (N678, N35_t13, N494_t2);
and AND2_47 (N681, N35_t14, N511_t2);
and AND2_48 (N684, N35_t15, N528_t2);
and AND2_49 (N687, N52_t0, N273_t3);
and AND2_50 (N690, N52_t1, N290_t3);
and AND2_51 (N693, N52_t2, N307_t3);
and AND2_52 (N696, N52_t3, N324_t3);
and AND2_53 (N699, N52_t4, N341_t3);
and AND2_54 (N702, N52_t5, N358_t3);
and AND2_55 (N705, N52_t6, N375_t3);
and AND2_56 (N708, N52_t7, N392_t3);
and AND2_57 (N711, N52_t8, N409_t3);
and AND2_58 (N714, N52_t9, N426_t3);
and AND2_59 (N717, N52_t10, N443_t3);
and AND2_60 (N720, N52_t11, N460_t3);
and AND2_61 (N723, N52_t12, N477_t3);
and AND2_62 (N726, N52_t13, N494_t3);
and AND2_63 (N729, N52_t14, N511_t3);
and AND2_64 (N732, N52_t15, N528_t3);
and AND2_65 (N735, N69_t0, N273_t4);
and AND2_66 (N738, N69_t1, N290_t4);
and AND2_67 (N741, N69_t2, N307_t4);
and AND2_68 (N744, N69_t3, N324_t4);
and AND2_69 (N747, N69_t4, N341_t4);
and AND2_70 (N750, N69_t5, N358_t4);
and AND2_71 (N753, N69_t6, N375_t4);
and AND2_72 (N756, N69_t7, N392_t4);
and AND2_73 (N759, N69_t8, N409_t4);
and AND2_74 (N762, N69_t9, N426_t4);
and AND2_75 (N765, N69_t10, N443_t4);
and AND2_76 (N768, N69_t11, N460_t4);
and AND2_77 (N771, N69_t12, N477_t4);
and AND2_78 (N774, N69_t13, N494_t4);
and AND2_79 (N777, N69_t14, N511_t4);
and AND2_80 (N780, N69_t15, N528_t4);
and AND2_81 (N783, N86_t0, N273_t5);
and AND2_82 (N786, N86_t1, N290_t5);
and AND2_83 (N789, N86_t2, N307_t5);
and AND2_84 (N792, N86_t3, N324_t5);
and AND2_85 (N795, N86_t4, N341_t5);
and AND2_86 (N798, N86_t5, N358_t5);
and AND2_87 (N801, N86_t6, N375_t5);
and AND2_88 (N804, N86_t7, N392_t5);
and AND2_89 (N807, N86_t8, N409_t5);
and AND2_90 (N810, N86_t9, N426_t5);
and AND2_91 (N813, N86_t10, N443_t5);
and AND2_92 (N816, N86_t11, N460_t5);
and AND2_93 (N819, N86_t12, N477_t5);
and AND2_94 (N822, N86_t13, N494_t5);
and AND2_95 (N825, N86_t14, N511_t5);
and AND2_96 (N828, N86_t15, N528_t5);
and AND2_97 (N831, N103_t0, N273_t6);
and AND2_98 (N834, N103_t1, N290_t6);
and AND2_99 (N837, N103_t2, N307_t6);
and AND2_100 (N840, N103_t3, N324_t6);
and AND2_101 (N843, N103_t4, N341_t6);
and AND2_102 (N846, N103_t5, N358_t6);
and AND2_103 (N849, N103_t6, N375_t6);
and AND2_104 (N852, N103_t7, N392_t6);
and AND2_105 (N855, N103_t8, N409_t6);
and AND2_106 (N858, N103_t9, N426_t6);
and AND2_107 (N861, N103_t10, N443_t6);
and AND2_108 (N864, N103_t11, N460_t6);
and AND2_109 (N867, N103_t12, N477_t6);
and AND2_110 (N870, N103_t13, N494_t6);
and AND2_111 (N873, N103_t14, N511_t6);
and AND2_112 (N876, N103_t15, N528_t6);
and AND2_113 (N879, N120_t0, N273_t7);
and AND2_114 (N882, N120_t1, N290_t7);
and AND2_115 (N885, N120_t2, N307_t7);
and AND2_116 (N888, N120_t3, N324_t7);
and AND2_117 (N891, N120_t4, N341_t7);
and AND2_118 (N894, N120_t5, N358_t7);
and AND2_119 (N897, N120_t6, N375_t7);
and AND2_120 (N900, N120_t7, N392_t7);
and AND2_121 (N903, N120_t8, N409_t7);
and AND2_122 (N906, N120_t9, N426_t7);
and AND2_123 (N909, N120_t10, N443_t7);
and AND2_124 (N912, N120_t11, N460_t7);
and AND2_125 (N915, N120_t12, N477_t7);
and AND2_126 (N918, N120_t13, N494_t7);
and AND2_127 (N921, N120_t14, N511_t7);
and AND2_128 (N924, N120_t15, N528_t7);
and AND2_129 (N927, N137_t0, N273_t8);
and AND2_130 (N930, N137_t1, N290_t8);
and AND2_131 (N933, N137_t2, N307_t8);
and AND2_132 (N936, N137_t3, N324_t8);
and AND2_133 (N939, N137_t4, N341_t8);
and AND2_134 (N942, N137_t5, N358_t8);
and AND2_135 (N945, N137_t6, N375_t8);
and AND2_136 (N948, N137_t7, N392_t8);
and AND2_137 (N951, N137_t8, N409_t8);
and AND2_138 (N954, N137_t9, N426_t8);
and AND2_139 (N957, N137_t10, N443_t8);
and AND2_140 (N960, N137_t11, N460_t8);
and AND2_141 (N963, N137_t12, N477_t8);
and AND2_142 (N966, N137_t13, N494_t8);
and AND2_143 (N969, N137_t14, N511_t8);
and AND2_144 (N972, N137_t15, N528_t8);
and AND2_145 (N975, N154_t0, N273_t9);
and AND2_146 (N978, N154_t1, N290_t9);
and AND2_147 (N981, N154_t2, N307_t9);
and AND2_148 (N984, N154_t3, N324_t9);
and AND2_149 (N987, N154_t4, N341_t9);
and AND2_150 (N990, N154_t5, N358_t9);
and AND2_151 (N993, N154_t6, N375_t9);
and AND2_152 (N996, N154_t7, N392_t9);
and AND2_153 (N999, N154_t8, N409_t9);
and AND2_154 (N1002, N154_t9, N426_t9);
and AND2_155 (N1005, N154_t10, N443_t9);
and AND2_156 (N1008, N154_t11, N460_t9);
and AND2_157 (N1011, N154_t12, N477_t9);
and AND2_158 (N1014, N154_t13, N494_t9);
and AND2_159 (N1017, N154_t14, N511_t9);
and AND2_160 (N1020, N154_t15, N528_t9);
and AND2_161 (N1023, N171_t0, N273_t10);
and AND2_162 (N1026, N171_t1, N290_t10);
and AND2_163 (N1029, N171_t2, N307_t10);
and AND2_164 (N1032, N171_t3, N324_t10);
and AND2_165 (N1035, N171_t4, N341_t10);
and AND2_166 (N1038, N171_t5, N358_t10);
and AND2_167 (N1041, N171_t6, N375_t10);
and AND2_168 (N1044, N171_t7, N392_t10);
and AND2_169 (N1047, N171_t8, N409_t10);
and AND2_170 (N1050, N171_t9, N426_t10);
and AND2_171 (N1053, N171_t10, N443_t10);
and AND2_172 (N1056, N171_t11, N460_t10);
and AND2_173 (N1059, N171_t12, N477_t10);
and AND2_174 (N1062, N171_t13, N494_t10);
and AND2_175 (N1065, N171_t14, N511_t10);
and AND2_176 (N1068, N171_t15, N528_t10);
and AND2_177 (N1071, N188_t0, N273_t11);
and AND2_178 (N1074, N188_t1, N290_t11);
and AND2_179 (N1077, N188_t2, N307_t11);
and AND2_180 (N1080, N188_t3, N324_t11);
and AND2_181 (N1083, N188_t4, N341_t11);
and AND2_182 (N1086, N188_t5, N358_t11);
and AND2_183 (N1089, N188_t6, N375_t11);
and AND2_184 (N1092, N188_t7, N392_t11);
and AND2_185 (N1095, N188_t8, N409_t11);
and AND2_186 (N1098, N188_t9, N426_t11);
and AND2_187 (N1101, N188_t10, N443_t11);
and AND2_188 (N1104, N188_t11, N460_t11);
and AND2_189 (N1107, N188_t12, N477_t11);
and AND2_190 (N1110, N188_t13, N494_t11);
and AND2_191 (N1113, N188_t14, N511_t11);
and AND2_192 (N1116, N188_t15, N528_t11);
and AND2_193 (N1119, N205_t0, N273_t12);
and AND2_194 (N1122, N205_t1, N290_t12);
and AND2_195 (N1125, N205_t2, N307_t12);
and AND2_196 (N1128, N205_t3, N324_t12);
and AND2_197 (N1131, N205_t4, N341_t12);
and AND2_198 (N1134, N205_t5, N358_t12);
and AND2_199 (N1137, N205_t6, N375_t12);
and AND2_200 (N1140, N205_t7, N392_t12);
and AND2_201 (N1143, N205_t8, N409_t12);
and AND2_202 (N1146, N205_t9, N426_t12);
and AND2_203 (N1149, N205_t10, N443_t12);
and AND2_204 (N1152, N205_t11, N460_t12);
and AND2_205 (N1155, N205_t12, N477_t12);
and AND2_206 (N1158, N205_t13, N494_t12);
and AND2_207 (N1161, N205_t14, N511_t12);
and AND2_208 (N1164, N205_t15, N528_t12);
and AND2_209 (N1167, N222_t0, N273_t13);
and AND2_210 (N1170, N222_t1, N290_t13);
and AND2_211 (N1173, N222_t2, N307_t13);
and AND2_212 (N1176, N222_t3, N324_t13);
and AND2_213 (N1179, N222_t4, N341_t13);
and AND2_214 (N1182, N222_t5, N358_t13);
and AND2_215 (N1185, N222_t6, N375_t13);
and AND2_216 (N1188, N222_t7, N392_t13);
and AND2_217 (N1191, N222_t8, N409_t13);
and AND2_218 (N1194, N222_t9, N426_t13);
and AND2_219 (N1197, N222_t10, N443_t13);
and AND2_220 (N1200, N222_t11, N460_t13);
and AND2_221 (N1203, N222_t12, N477_t13);
and AND2_222 (N1206, N222_t13, N494_t13);
and AND2_223 (N1209, N222_t14, N511_t13);
and AND2_224 (N1212, N222_t15, N528_t13);
and AND2_225 (N1215, N239_t0, N273_t14);
and AND2_226 (N1218, N239_t1, N290_t14);
and AND2_227 (N1221, N239_t2, N307_t14);
and AND2_228 (N1224, N239_t3, N324_t14);
and AND2_229 (N1227, N239_t4, N341_t14);
and AND2_230 (N1230, N239_t5, N358_t14);
and AND2_231 (N1233, N239_t6, N375_t14);
and AND2_232 (N1236, N239_t7, N392_t14);
and AND2_233 (N1239, N239_t8, N409_t14);
and AND2_234 (N1242, N239_t9, N426_t14);
and AND2_235 (N1245, N239_t10, N443_t14);
and AND2_236 (N1248, N239_t11, N460_t14);
and AND2_237 (N1251, N239_t12, N477_t14);
and AND2_238 (N1254, N239_t13, N494_t14);
and AND2_239 (N1257, N239_t14, N511_t14);
and AND2_240 (N1260, N239_t15, N528_t14);
and AND2_241 (N1263, N256_t0, N273_t15);
and AND2_242 (N1266, N256_t1, N290_t15);
and AND2_243 (N1269, N256_t2, N307_t15);
and AND2_244 (N1272, N256_t3, N324_t15);
and AND2_245 (N1275, N256_t4, N341_t15);
and AND2_246 (N1278, N256_t5, N358_t15);
and AND2_247 (N1281, N256_t6, N375_t15);
and AND2_248 (N1284, N256_t7, N392_t15);
and AND2_249 (N1287, N256_t8, N409_t15);
and AND2_250 (N1290, N256_t9, N426_t15);
and AND2_251 (N1293, N256_t10, N443_t15);
and AND2_252 (N1296, N256_t11, N460_t15);
and AND2_253 (N1299, N256_t12, N477_t15);
and AND2_254 (N1302, N256_t13, N494_t15);
and AND2_255 (N1305, N256_t14, N511_t15);
and AND2_256 (N1308, N256_t15, N528_t15);
not NOT1_257 (N1311, N591_t0);
not NOT1_258 (N1315, N639_t0);
not NOT1_259 (N1319, N687_t0);
not NOT1_260 (N1323, N735_t0);
not NOT1_261 (N1327, N783_t0);
not NOT1_262 (N1331, N831_t0);
not NOT1_263 (N1335, N879_t0);
not NOT1_264 (N1339, N927_t0);
not NOT1_265 (N1343, N975_t0);
not NOT1_266 (N1347, N1023_t0);
not NOT1_267 (N1351, N1071_t0);
not NOT1_268 (N1355, N1119_t0);
not NOT1_269 (N1359, N1167_t0);
not NOT1_270 (N1363, N1215_t0);
not NOT1_271 (N1367, N1263_t0);
nor NOR2_272 (N1371, N591_t1, N1311_t0);
not NOT1_273 (N1372, N1311_t1);
nor NOR2_274 (N1373, N639_t1, N1315_t0);
not NOT1_275 (N1374, N1315_t1);
nor NOR2_276 (N1375, N687_t1, N1319_t0);
not NOT1_277 (N1376, N1319_t1);
nor NOR2_278 (N1377, N735_t1, N1323_t0);
not NOT1_279 (N1378, N1323_t1);
nor NOR2_280 (N1379, N783_t1, N1327_t0);
not NOT1_281 (N1380, N1327_t1);
nor NOR2_282 (N1381, N831_t1, N1331_t0);
not NOT1_283 (N1382, N1331_t1);
nor NOR2_284 (N1383, N879_t1, N1335_t0);
not NOT1_285 (N1384, N1335_t1);
nor NOR2_286 (N1385, N927_t1, N1339_t0);
not NOT1_287 (N1386, N1339_t1);
nor NOR2_288 (N1387, N975_t1, N1343_t0);
not NOT1_289 (N1388, N1343_t1);
nor NOR2_290 (N1389, N1023_t1, N1347_t0);
not NOT1_291 (N1390, N1347_t1);
nor NOR2_292 (N1391, N1071_t1, N1351_t0);
not NOT1_293 (N1392, N1351_t1);
nor NOR2_294 (N1393, N1119_t1, N1355_t0);
not NOT1_295 (N1394, N1355_t1);
nor NOR2_296 (N1395, N1167_t1, N1359_t0);
not NOT1_297 (N1396, N1359_t1);
nor NOR2_298 (N1397, N1215_t1, N1363_t0);
not NOT1_299 (N1398, N1363_t1);
nor NOR2_300 (N1399, N1263_t1, N1367_t0);
not NOT1_301 (N1400, N1367_t1);
nor NOR2_302 (N1401, N1371, N1372);
nor NOR2_303 (N1404, N1373, N1374);
nor NOR2_304 (N1407, N1375, N1376);
nor NOR2_305 (N1410, N1377, N1378);
nor NOR2_306 (N1413, N1379, N1380);
nor NOR2_307 (N1416, N1381, N1382);
nor NOR2_308 (N1419, N1383, N1384);
nor NOR2_309 (N1422, N1385, N1386);
nor NOR2_310 (N1425, N1387, N1388);
nor NOR2_311 (N1428, N1389, N1390);
nor NOR2_312 (N1431, N1391, N1392);
nor NOR2_313 (N1434, N1393, N1394);
nor NOR2_314 (N1437, N1395, N1396);
nor NOR2_315 (N1440, N1397, N1398);
nor NOR2_316 (N1443, N1399, N1400);
nor NOR2_317 (N1446, N1401_t0, N546_t0);
nor NOR2_318 (N1450, N1404_t0, N594_t0);
nor NOR2_319 (N1454, N1407_t0, N642_t0);
nor NOR2_320 (N1458, N1410_t0, N690_t0);
nor NOR2_321 (N1462, N1413_t0, N738_t0);
nor NOR2_322 (N1466, N1416_t0, N786_t0);
nor NOR2_323 (N1470, N1419_t0, N834_t0);
nor NOR2_324 (N1474, N1422_t0, N882_t0);
nor NOR2_325 (N1478, N1425_t0, N930_t0);
nor NOR2_326 (N1482, N1428_t0, N978_t0);
nor NOR2_327 (N1486, N1431_t0, N1026_t0);
nor NOR2_328 (N1490, N1434_t0, N1074_t0);
nor NOR2_329 (N1494, N1437_t0, N1122_t0);
nor NOR2_330 (N1498, N1440_t0, N1170_t0);
nor NOR2_331 (N1502, N1443_t0, N1218_t0);
nor NOR2_332 (N1506, N1401_t1, N1446_t0);
nor NOR2_333 (N1507, N1446_t1, N546_t1);
nor NOR2_334 (N1508, N1311_t2, N1446_t2);
nor NOR2_335 (N1511, N1404_t1, N1450_t0);
nor NOR2_336 (N1512, N1450_t1, N594_t1);
nor NOR2_337 (N1513, N1315_t2, N1450_t2);
nor NOR2_338 (N1516, N1407_t1, N1454_t0);
nor NOR2_339 (N1517, N1454_t1, N642_t1);
nor NOR2_340 (N1518, N1319_t2, N1454_t2);
nor NOR2_341 (N1521, N1410_t1, N1458_t0);
nor NOR2_342 (N1522, N1458_t1, N690_t1);
nor NOR2_343 (N1523, N1323_t2, N1458_t2);
nor NOR2_344 (N1526, N1413_t1, N1462_t0);
nor NOR2_345 (N1527, N1462_t1, N738_t1);
nor NOR2_346 (N1528, N1327_t2, N1462_t2);
nor NOR2_347 (N1531, N1416_t1, N1466_t0);
nor NOR2_348 (N1532, N1466_t1, N786_t1);
nor NOR2_349 (N1533, N1331_t2, N1466_t2);
nor NOR2_350 (N1536, N1419_t1, N1470_t0);
nor NOR2_351 (N1537, N1470_t1, N834_t1);
nor NOR2_352 (N1538, N1335_t2, N1470_t2);
nor NOR2_353 (N1541, N1422_t1, N1474_t0);
nor NOR2_354 (N1542, N1474_t1, N882_t1);
nor NOR2_355 (N1543, N1339_t2, N1474_t2);
nor NOR2_356 (N1546, N1425_t1, N1478_t0);
nor NOR2_357 (N1547, N1478_t1, N930_t1);
nor NOR2_358 (N1548, N1343_t2, N1478_t2);
nor NOR2_359 (N1551, N1428_t1, N1482_t0);
nor NOR2_360 (N1552, N1482_t1, N978_t1);
nor NOR2_361 (N1553, N1347_t2, N1482_t2);
nor NOR2_362 (N1556, N1431_t1, N1486_t0);
nor NOR2_363 (N1557, N1486_t1, N1026_t1);
nor NOR2_364 (N1558, N1351_t2, N1486_t2);
nor NOR2_365 (N1561, N1434_t1, N1490_t0);
nor NOR2_366 (N1562, N1490_t1, N1074_t1);
nor NOR2_367 (N1563, N1355_t2, N1490_t2);
nor NOR2_368 (N1566, N1437_t1, N1494_t0);
nor NOR2_369 (N1567, N1494_t1, N1122_t1);
nor NOR2_370 (N1568, N1359_t2, N1494_t2);
nor NOR2_371 (N1571, N1440_t1, N1498_t0);
nor NOR2_372 (N1572, N1498_t1, N1170_t1);
nor NOR2_373 (N1573, N1363_t2, N1498_t2);
nor NOR2_374 (N1576, N1443_t1, N1502_t0);
nor NOR2_375 (N1577, N1502_t1, N1218_t1);
nor NOR2_376 (N1578, N1367_t2, N1502_t2);
nor NOR2_377 (N1581, N1506, N1507);
nor NOR2_378 (N1582, N1511, N1512);
nor NOR2_379 (N1585, N1516, N1517);
nor NOR2_380 (N1588, N1521, N1522);
nor NOR2_381 (N1591, N1526, N1527);
nor NOR2_382 (N1594, N1531, N1532);
nor NOR2_383 (N1597, N1536, N1537);
nor NOR2_384 (N1600, N1541, N1542);
nor NOR2_385 (N1603, N1546, N1547);
nor NOR2_386 (N1606, N1551, N1552);
nor NOR2_387 (N1609, N1556, N1557);
nor NOR2_388 (N1612, N1561, N1562);
nor NOR2_389 (N1615, N1566, N1567);
nor NOR2_390 (N1618, N1571, N1572);
nor NOR2_391 (N1621, N1576, N1577);
nor NOR2_392 (N1624, N1266_t0, N1578_t0);
nor NOR2_393 (N1628, N1582_t0, N1508_t0);
nor NOR2_394 (N1632, N1585_t0, N1513_t0);
nor NOR2_395 (N1636, N1588_t0, N1518_t0);
nor NOR2_396 (N1640, N1591_t0, N1523_t0);
nor NOR2_397 (N1644, N1594_t0, N1528_t0);
nor NOR2_398 (N1648, N1597_t0, N1533_t0);
nor NOR2_399 (N1652, N1600_t0, N1538_t0);
nor NOR2_400 (N1656, N1603_t0, N1543_t0);
nor NOR2_401 (N1660, N1606_t0, N1548_t0);
nor NOR2_402 (N1664, N1609_t0, N1553_t0);
nor NOR2_403 (N1668, N1612_t0, N1558_t0);
nor NOR2_404 (N1672, N1615_t0, N1563_t0);
nor NOR2_405 (N1676, N1618_t0, N1568_t0);
nor NOR2_406 (N1680, N1621_t0, N1573_t0);
nor NOR2_407 (N1684, N1266_t1, N1624_t0);
nor NOR2_408 (N1685, N1624_t1, N1578_t1);
nor NOR2_409 (N1686, N1582_t1, N1628_t0);
nor NOR2_410 (N1687, N1628_t1, N1508_t1);
nor NOR2_411 (N1688, N1585_t1, N1632_t0);
nor NOR2_412 (N1689, N1632_t1, N1513_t1);
nor NOR2_413 (N1690, N1588_t1, N1636_t0);
nor NOR2_414 (N1691, N1636_t1, N1518_t1);
nor NOR2_415 (N1692, N1591_t1, N1640_t0);
nor NOR2_416 (N1693, N1640_t1, N1523_t1);
nor NOR2_417 (N1694, N1594_t1, N1644_t0);
nor NOR2_418 (N1695, N1644_t1, N1528_t1);
nor NOR2_419 (N1696, N1597_t1, N1648_t0);
nor NOR2_420 (N1697, N1648_t1, N1533_t1);
nor NOR2_421 (N1698, N1600_t1, N1652_t0);
nor NOR2_422 (N1699, N1652_t1, N1538_t1);
nor NOR2_423 (N1700, N1603_t1, N1656_t0);
nor NOR2_424 (N1701, N1656_t1, N1543_t1);
nor NOR2_425 (N1702, N1606_t1, N1660_t0);
nor NOR2_426 (N1703, N1660_t1, N1548_t1);
nor NOR2_427 (N1704, N1609_t1, N1664_t0);
nor NOR2_428 (N1705, N1664_t1, N1553_t1);
nor NOR2_429 (N1706, N1612_t1, N1668_t0);
nor NOR2_430 (N1707, N1668_t1, N1558_t1);
nor NOR2_431 (N1708, N1615_t1, N1672_t0);
nor NOR2_432 (N1709, N1672_t1, N1563_t1);
nor NOR2_433 (N1710, N1618_t1, N1676_t0);
nor NOR2_434 (N1711, N1676_t1, N1568_t1);
nor NOR2_435 (N1712, N1621_t1, N1680_t0);
nor NOR2_436 (N1713, N1680_t1, N1573_t1);
nor NOR2_437 (N1714, N1684, N1685);
nor NOR2_438 (N1717, N1686, N1687);
nor NOR2_439 (N1720, N1688, N1689);
nor NOR2_440 (N1723, N1690, N1691);
nor NOR2_441 (N1726, N1692, N1693);
nor NOR2_442 (N1729, N1694, N1695);
nor NOR2_443 (N1732, N1696, N1697);
nor NOR2_444 (N1735, N1698, N1699);
nor NOR2_445 (N1738, N1700, N1701);
nor NOR2_446 (N1741, N1702, N1703);
nor NOR2_447 (N1744, N1704, N1705);
nor NOR2_448 (N1747, N1706, N1707);
nor NOR2_449 (N1750, N1708, N1709);
nor NOR2_450 (N1753, N1710, N1711);
nor NOR2_451 (N1756, N1712, N1713);
nor NOR2_452 (N1759, N1714_t0, N1221_t0);
nor NOR2_453 (N1763, N1717_t0, N549_t0);
nor NOR2_454 (N1767, N1720_t0, N597_t0);
nor NOR2_455 (N1771, N1723_t0, N645_t0);
nor NOR2_456 (N1775, N1726_t0, N693_t0);
nor NOR2_457 (N1779, N1729_t0, N741_t0);
nor NOR2_458 (N1783, N1732_t0, N789_t0);
nor NOR2_459 (N1787, N1735_t0, N837_t0);
nor NOR2_460 (N1791, N1738_t0, N885_t0);
nor NOR2_461 (N1795, N1741_t0, N933_t0);
nor NOR2_462 (N1799, N1744_t0, N981_t0);
nor NOR2_463 (N1803, N1747_t0, N1029_t0);
nor NOR2_464 (N1807, N1750_t0, N1077_t0);
nor NOR2_465 (N1811, N1753_t0, N1125_t0);
nor NOR2_466 (N1815, N1756_t0, N1173_t0);
nor NOR2_467 (N1819, N1714_t1, N1759_t0);
nor NOR2_468 (N1820, N1759_t1, N1221_t1);
nor NOR2_469 (N1821, N1624_t2, N1759_t2);
nor NOR2_470 (N1824, N1717_t1, N1763_t0);
nor NOR2_471 (N1825, N1763_t1, N549_t1);
nor NOR2_472 (N1826, N1628_t2, N1763_t2);
nor NOR2_473 (N1829, N1720_t1, N1767_t0);
nor NOR2_474 (N1830, N1767_t1, N597_t1);
nor NOR2_475 (N1831, N1632_t2, N1767_t2);
nor NOR2_476 (N1834, N1723_t1, N1771_t0);
nor NOR2_477 (N1835, N1771_t1, N645_t1);
nor NOR2_478 (N1836, N1636_t2, N1771_t2);
nor NOR2_479 (N1839, N1726_t1, N1775_t0);
nor NOR2_480 (N1840, N1775_t1, N693_t1);
nor NOR2_481 (N1841, N1640_t2, N1775_t2);
nor NOR2_482 (N1844, N1729_t1, N1779_t0);
nor NOR2_483 (N1845, N1779_t1, N741_t1);
nor NOR2_484 (N1846, N1644_t2, N1779_t2);
nor NOR2_485 (N1849, N1732_t1, N1783_t0);
nor NOR2_486 (N1850, N1783_t1, N789_t1);
nor NOR2_487 (N1851, N1648_t2, N1783_t2);
nor NOR2_488 (N1854, N1735_t1, N1787_t0);
nor NOR2_489 (N1855, N1787_t1, N837_t1);
nor NOR2_490 (N1856, N1652_t2, N1787_t2);
nor NOR2_491 (N1859, N1738_t1, N1791_t0);
nor NOR2_492 (N1860, N1791_t1, N885_t1);
nor NOR2_493 (N1861, N1656_t2, N1791_t2);
nor NOR2_494 (N1864, N1741_t1, N1795_t0);
nor NOR2_495 (N1865, N1795_t1, N933_t1);
nor NOR2_496 (N1866, N1660_t2, N1795_t2);
nor NOR2_497 (N1869, N1744_t1, N1799_t0);
nor NOR2_498 (N1870, N1799_t1, N981_t1);
nor NOR2_499 (N1871, N1664_t2, N1799_t2);
nor NOR2_500 (N1874, N1747_t1, N1803_t0);
nor NOR2_501 (N1875, N1803_t1, N1029_t1);
nor NOR2_502 (N1876, N1668_t2, N1803_t2);
nor NOR2_503 (N1879, N1750_t1, N1807_t0);
nor NOR2_504 (N1880, N1807_t1, N1077_t1);
nor NOR2_505 (N1881, N1672_t2, N1807_t2);
nor NOR2_506 (N1884, N1753_t1, N1811_t0);
nor NOR2_507 (N1885, N1811_t1, N1125_t1);
nor NOR2_508 (N1886, N1676_t2, N1811_t2);
nor NOR2_509 (N1889, N1756_t1, N1815_t0);
nor NOR2_510 (N1890, N1815_t1, N1173_t1);
nor NOR2_511 (N1891, N1680_t2, N1815_t2);
nor NOR2_512 (N1894, N1819, N1820);
nor NOR2_513 (N1897, N1269_t0, N1821_t0);
nor NOR2_514 (N1901, N1824, N1825);
nor NOR2_515 (N1902, N1829, N1830);
nor NOR2_516 (N1905, N1834, N1835);
nor NOR2_517 (N1908, N1839, N1840);
nor NOR2_518 (N1911, N1844, N1845);
nor NOR2_519 (N1914, N1849, N1850);
nor NOR2_520 (N1917, N1854, N1855);
nor NOR2_521 (N1920, N1859, N1860);
nor NOR2_522 (N1923, N1864, N1865);
nor NOR2_523 (N1926, N1869, N1870);
nor NOR2_524 (N1929, N1874, N1875);
nor NOR2_525 (N1932, N1879, N1880);
nor NOR2_526 (N1935, N1884, N1885);
nor NOR2_527 (N1938, N1889, N1890);
nor NOR2_528 (N1941, N1894_t0, N1891_t0);
nor NOR2_529 (N1945, N1269_t1, N1897_t0);
nor NOR2_530 (N1946, N1897_t1, N1821_t1);
nor NOR2_531 (N1947, N1902_t0, N1826_t0);
nor NOR2_532 (N1951, N1905_t0, N1831_t0);
nor NOR2_533 (N1955, N1908_t0, N1836_t0);
nor NOR2_534 (N1959, N1911_t0, N1841_t0);
nor NOR2_535 (N1963, N1914_t0, N1846_t0);
nor NOR2_536 (N1967, N1917_t0, N1851_t0);
nor NOR2_537 (N1971, N1920_t0, N1856_t0);
nor NOR2_538 (N1975, N1923_t0, N1861_t0);
nor NOR2_539 (N1979, N1926_t0, N1866_t0);
nor NOR2_540 (N1983, N1929_t0, N1871_t0);
nor NOR2_541 (N1987, N1932_t0, N1876_t0);
nor NOR2_542 (N1991, N1935_t0, N1881_t0);
nor NOR2_543 (N1995, N1938_t0, N1886_t0);
nor NOR2_544 (N1999, N1894_t1, N1941_t0);
nor NOR2_545 (N2000, N1941_t1, N1891_t1);
nor NOR2_546 (N2001, N1945, N1946);
nor NOR2_547 (N2004, N1902_t1, N1947_t0);
nor NOR2_548 (N2005, N1947_t1, N1826_t1);
nor NOR2_549 (N2006, N1905_t1, N1951_t0);
nor NOR2_550 (N2007, N1951_t1, N1831_t1);
nor NOR2_551 (N2008, N1908_t1, N1955_t0);
nor NOR2_552 (N2009, N1955_t1, N1836_t1);
nor NOR2_553 (N2010, N1911_t1, N1959_t0);
nor NOR2_554 (N2011, N1959_t1, N1841_t1);
nor NOR2_555 (N2012, N1914_t1, N1963_t0);
nor NOR2_556 (N2013, N1963_t1, N1846_t1);
nor NOR2_557 (N2014, N1917_t1, N1967_t0);
nor NOR2_558 (N2015, N1967_t1, N1851_t1);
nor NOR2_559 (N2016, N1920_t1, N1971_t0);
nor NOR2_560 (N2017, N1971_t1, N1856_t1);
nor NOR2_561 (N2018, N1923_t1, N1975_t0);
nor NOR2_562 (N2019, N1975_t1, N1861_t1);
nor NOR2_563 (N2020, N1926_t1, N1979_t0);
nor NOR2_564 (N2021, N1979_t1, N1866_t1);
nor NOR2_565 (N2022, N1929_t1, N1983_t0);
nor NOR2_566 (N2023, N1983_t1, N1871_t1);
nor NOR2_567 (N2024, N1932_t1, N1987_t0);
nor NOR2_568 (N2025, N1987_t1, N1876_t1);
nor NOR2_569 (N2026, N1935_t1, N1991_t0);
nor NOR2_570 (N2027, N1991_t1, N1881_t1);
nor NOR2_571 (N2028, N1938_t1, N1995_t0);
nor NOR2_572 (N2029, N1995_t1, N1886_t1);
nor NOR2_573 (N2030, N1999, N2000);
nor NOR2_574 (N2033, N2001_t0, N1224_t0);
nor NOR2_575 (N2037, N2004, N2005);
nor NOR2_576 (N2040, N2006, N2007);
nor NOR2_577 (N2043, N2008, N2009);
nor NOR2_578 (N2046, N2010, N2011);
nor NOR2_579 (N2049, N2012, N2013);
nor NOR2_580 (N2052, N2014, N2015);
nor NOR2_581 (N2055, N2016, N2017);
nor NOR2_582 (N2058, N2018, N2019);
nor NOR2_583 (N2061, N2020, N2021);
nor NOR2_584 (N2064, N2022, N2023);
nor NOR2_585 (N2067, N2024, N2025);
nor NOR2_586 (N2070, N2026, N2027);
nor NOR2_587 (N2073, N2028, N2029);
nor NOR2_588 (N2076, N2030_t0, N1176_t0);
nor NOR2_589 (N2080, N2001_t1, N2033_t0);
nor NOR2_590 (N2081, N2033_t1, N1224_t1);
nor NOR2_591 (N2082, N1897_t2, N2033_t2);
nor NOR2_592 (N2085, N2037_t0, N552_t0);
nor NOR2_593 (N2089, N2040_t0, N600_t0);
nor NOR2_594 (N2093, N2043_t0, N648_t0);
nor NOR2_595 (N2097, N2046_t0, N696_t0);
nor NOR2_596 (N2101, N2049_t0, N744_t0);
nor NOR2_597 (N2105, N2052_t0, N792_t0);
nor NOR2_598 (N2109, N2055_t0, N840_t0);
nor NOR2_599 (N2113, N2058_t0, N888_t0);
nor NOR2_600 (N2117, N2061_t0, N936_t0);
nor NOR2_601 (N2121, N2064_t0, N984_t0);
nor NOR2_602 (N2125, N2067_t0, N1032_t0);
nor NOR2_603 (N2129, N2070_t0, N1080_t0);
nor NOR2_604 (N2133, N2073_t0, N1128_t0);
nor NOR2_605 (N2137, N2030_t1, N2076_t0);
nor NOR2_606 (N2138, N2076_t1, N1176_t1);
nor NOR2_607 (N2139, N1941_t2, N2076_t2);
nor NOR2_608 (N2142, N2080, N2081);
nor NOR2_609 (N2145, N1272_t0, N2082_t0);
nor NOR2_610 (N2149, N2037_t1, N2085_t0);
nor NOR2_611 (N2150, N2085_t1, N552_t1);
nor NOR2_612 (N2151, N1947_t2, N2085_t2);
nor NOR2_613 (N2154, N2040_t1, N2089_t0);
nor NOR2_614 (N2155, N2089_t1, N600_t1);
nor NOR2_615 (N2156, N1951_t2, N2089_t2);
nor NOR2_616 (N2159, N2043_t1, N2093_t0);
nor NOR2_617 (N2160, N2093_t1, N648_t1);
nor NOR2_618 (N2161, N1955_t2, N2093_t2);
nor NOR2_619 (N2164, N2046_t1, N2097_t0);
nor NOR2_620 (N2165, N2097_t1, N696_t1);
nor NOR2_621 (N2166, N1959_t2, N2097_t2);
nor NOR2_622 (N2169, N2049_t1, N2101_t0);
nor NOR2_623 (N2170, N2101_t1, N744_t1);
nor NOR2_624 (N2171, N1963_t2, N2101_t2);
nor NOR2_625 (N2174, N2052_t1, N2105_t0);
nor NOR2_626 (N2175, N2105_t1, N792_t1);
nor NOR2_627 (N2176, N1967_t2, N2105_t2);
nor NOR2_628 (N2179, N2055_t1, N2109_t0);
nor NOR2_629 (N2180, N2109_t1, N840_t1);
nor NOR2_630 (N2181, N1971_t2, N2109_t2);
nor NOR2_631 (N2184, N2058_t1, N2113_t0);
nor NOR2_632 (N2185, N2113_t1, N888_t1);
nor NOR2_633 (N2186, N1975_t2, N2113_t2);
nor NOR2_634 (N2189, N2061_t1, N2117_t0);
nor NOR2_635 (N2190, N2117_t1, N936_t1);
nor NOR2_636 (N2191, N1979_t2, N2117_t2);
nor NOR2_637 (N2194, N2064_t1, N2121_t0);
nor NOR2_638 (N2195, N2121_t1, N984_t1);
nor NOR2_639 (N2196, N1983_t2, N2121_t2);
nor NOR2_640 (N2199, N2067_t1, N2125_t0);
nor NOR2_641 (N2200, N2125_t1, N1032_t1);
nor NOR2_642 (N2201, N1987_t2, N2125_t2);
nor NOR2_643 (N2204, N2070_t1, N2129_t0);
nor NOR2_644 (N2205, N2129_t1, N1080_t1);
nor NOR2_645 (N2206, N1991_t2, N2129_t2);
nor NOR2_646 (N2209, N2073_t1, N2133_t0);
nor NOR2_647 (N2210, N2133_t1, N1128_t1);
nor NOR2_648 (N2211, N1995_t2, N2133_t2);
nor NOR2_649 (N2214, N2137, N2138);
nor NOR2_650 (N2217, N2142_t0, N2139_t0);
nor NOR2_651 (N2221, N1272_t1, N2145_t0);
nor NOR2_652 (N2222, N2145_t1, N2082_t1);
nor NOR2_653 (N2223, N2149, N2150);
nor NOR2_654 (N2224, N2154, N2155);
nor NOR2_655 (N2227, N2159, N2160);
nor NOR2_656 (N2230, N2164, N2165);
nor NOR2_657 (N2233, N2169, N2170);
nor NOR2_658 (N2236, N2174, N2175);
nor NOR2_659 (N2239, N2179, N2180);
nor NOR2_660 (N2242, N2184, N2185);
nor NOR2_661 (N2245, N2189, N2190);
nor NOR2_662 (N2248, N2194, N2195);
nor NOR2_663 (N2251, N2199, N2200);
nor NOR2_664 (N2254, N2204, N2205);
nor NOR2_665 (N2257, N2209, N2210);
nor NOR2_666 (N2260, N2214_t0, N2211_t0);
nor NOR2_667 (N2264, N2142_t1, N2217_t0);
nor NOR2_668 (N2265, N2217_t1, N2139_t1);
nor NOR2_669 (N2266, N2221, N2222);
nor NOR2_670 (N2269, N2224_t0, N2151_t0);
nor NOR2_671 (N2273, N2227_t0, N2156_t0);
nor NOR2_672 (N2277, N2230_t0, N2161_t0);
nor NOR2_673 (N2281, N2233_t0, N2166_t0);
nor NOR2_674 (N2285, N2236_t0, N2171_t0);
nor NOR2_675 (N2289, N2239_t0, N2176_t0);
nor NOR2_676 (N2293, N2242_t0, N2181_t0);
nor NOR2_677 (N2297, N2245_t0, N2186_t0);
nor NOR2_678 (N2301, N2248_t0, N2191_t0);
nor NOR2_679 (N2305, N2251_t0, N2196_t0);
nor NOR2_680 (N2309, N2254_t0, N2201_t0);
nor NOR2_681 (N2313, N2257_t0, N2206_t0);
nor NOR2_682 (N2317, N2214_t1, N2260_t0);
nor NOR2_683 (N2318, N2260_t1, N2211_t1);
nor NOR2_684 (N2319, N2264, N2265);
nor NOR2_685 (N2322, N2266_t0, N1227_t0);
nor NOR2_686 (N2326, N2224_t1, N2269_t0);
nor NOR2_687 (N2327, N2269_t1, N2151_t1);
nor NOR2_688 (N2328, N2227_t1, N2273_t0);
nor NOR2_689 (N2329, N2273_t1, N2156_t1);
nor NOR2_690 (N2330, N2230_t1, N2277_t0);
nor NOR2_691 (N2331, N2277_t1, N2161_t1);
nor NOR2_692 (N2332, N2233_t1, N2281_t0);
nor NOR2_693 (N2333, N2281_t1, N2166_t1);
nor NOR2_694 (N2334, N2236_t1, N2285_t0);
nor NOR2_695 (N2335, N2285_t1, N2171_t1);
nor NOR2_696 (N2336, N2239_t1, N2289_t0);
nor NOR2_697 (N2337, N2289_t1, N2176_t1);
nor NOR2_698 (N2338, N2242_t1, N2293_t0);
nor NOR2_699 (N2339, N2293_t1, N2181_t1);
nor NOR2_700 (N2340, N2245_t1, N2297_t0);
nor NOR2_701 (N2341, N2297_t1, N2186_t1);
nor NOR2_702 (N2342, N2248_t1, N2301_t0);
nor NOR2_703 (N2343, N2301_t1, N2191_t1);
nor NOR2_704 (N2344, N2251_t1, N2305_t0);
nor NOR2_705 (N2345, N2305_t1, N2196_t1);
nor NOR2_706 (N2346, N2254_t1, N2309_t0);
nor NOR2_707 (N2347, N2309_t1, N2201_t1);
nor NOR2_708 (N2348, N2257_t1, N2313_t0);
nor NOR2_709 (N2349, N2313_t1, N2206_t1);
nor NOR2_710 (N2350, N2317, N2318);
nor NOR2_711 (N2353, N2319_t0, N1179_t0);
nor NOR2_712 (N2357, N2266_t1, N2322_t0);
nor NOR2_713 (N2358, N2322_t1, N1227_t1);
nor NOR2_714 (N2359, N2145_t2, N2322_t2);
nor NOR2_715 (N2362, N2326, N2327);
nor NOR2_716 (N2365, N2328, N2329);
nor NOR2_717 (N2368, N2330, N2331);
nor NOR2_718 (N2371, N2332, N2333);
nor NOR2_719 (N2374, N2334, N2335);
nor NOR2_720 (N2377, N2336, N2337);
nor NOR2_721 (N2380, N2338, N2339);
nor NOR2_722 (N2383, N2340, N2341);
nor NOR2_723 (N2386, N2342, N2343);
nor NOR2_724 (N2389, N2344, N2345);
nor NOR2_725 (N2392, N2346, N2347);
nor NOR2_726 (N2395, N2348, N2349);
nor NOR2_727 (N2398, N2350_t0, N1131_t0);
nor NOR2_728 (N2402, N2319_t1, N2353_t0);
nor NOR2_729 (N2403, N2353_t1, N1179_t1);
nor NOR2_730 (N2404, N2217_t2, N2353_t2);
nor NOR2_731 (N2407, N2357, N2358);
nor NOR2_732 (N2410, N1275_t0, N2359_t0);
nor NOR2_733 (N2414, N2362_t0, N555_t0);
nor NOR2_734 (N2418, N2365_t0, N603_t0);
nor NOR2_735 (N2422, N2368_t0, N651_t0);
nor NOR2_736 (N2426, N2371_t0, N699_t0);
nor NOR2_737 (N2430, N2374_t0, N747_t0);
nor NOR2_738 (N2434, N2377_t0, N795_t0);
nor NOR2_739 (N2438, N2380_t0, N843_t0);
nor NOR2_740 (N2442, N2383_t0, N891_t0);
nor NOR2_741 (N2446, N2386_t0, N939_t0);
nor NOR2_742 (N2450, N2389_t0, N987_t0);
nor NOR2_743 (N2454, N2392_t0, N1035_t0);
nor NOR2_744 (N2458, N2395_t0, N1083_t0);
nor NOR2_745 (N2462, N2350_t1, N2398_t0);
nor NOR2_746 (N2463, N2398_t1, N1131_t1);
nor NOR2_747 (N2464, N2260_t2, N2398_t2);
nor NOR2_748 (N2467, N2402, N2403);
nor NOR2_749 (N2470, N2407_t0, N2404_t0);
nor NOR2_750 (N2474, N1275_t1, N2410_t0);
nor NOR2_751 (N2475, N2410_t1, N2359_t1);
nor NOR2_752 (N2476, N2362_t1, N2414_t0);
nor NOR2_753 (N2477, N2414_t1, N555_t1);
nor NOR2_754 (N2478, N2269_t2, N2414_t2);
nor NOR2_755 (N2481, N2365_t1, N2418_t0);
nor NOR2_756 (N2482, N2418_t1, N603_t1);
nor NOR2_757 (N2483, N2273_t2, N2418_t2);
nor NOR2_758 (N2486, N2368_t1, N2422_t0);
nor NOR2_759 (N2487, N2422_t1, N651_t1);
nor NOR2_760 (N2488, N2277_t2, N2422_t2);
nor NOR2_761 (N2491, N2371_t1, N2426_t0);
nor NOR2_762 (N2492, N2426_t1, N699_t1);
nor NOR2_763 (N2493, N2281_t2, N2426_t2);
nor NOR2_764 (N2496, N2374_t1, N2430_t0);
nor NOR2_765 (N2497, N2430_t1, N747_t1);
nor NOR2_766 (N2498, N2285_t2, N2430_t2);
nor NOR2_767 (N2501, N2377_t1, N2434_t0);
nor NOR2_768 (N2502, N2434_t1, N795_t1);
nor NOR2_769 (N2503, N2289_t2, N2434_t2);
nor NOR2_770 (N2506, N2380_t1, N2438_t0);
nor NOR2_771 (N2507, N2438_t1, N843_t1);
nor NOR2_772 (N2508, N2293_t2, N2438_t2);
nor NOR2_773 (N2511, N2383_t1, N2442_t0);
nor NOR2_774 (N2512, N2442_t1, N891_t1);
nor NOR2_775 (N2513, N2297_t2, N2442_t2);
nor NOR2_776 (N2516, N2386_t1, N2446_t0);
nor NOR2_777 (N2517, N2446_t1, N939_t1);
nor NOR2_778 (N2518, N2301_t2, N2446_t2);
nor NOR2_779 (N2521, N2389_t1, N2450_t0);
nor NOR2_780 (N2522, N2450_t1, N987_t1);
nor NOR2_781 (N2523, N2305_t2, N2450_t2);
nor NOR2_782 (N2526, N2392_t1, N2454_t0);
nor NOR2_783 (N2527, N2454_t1, N1035_t1);
nor NOR2_784 (N2528, N2309_t2, N2454_t2);
nor NOR2_785 (N2531, N2395_t1, N2458_t0);
nor NOR2_786 (N2532, N2458_t1, N1083_t1);
nor NOR2_787 (N2533, N2313_t2, N2458_t2);
nor NOR2_788 (N2536, N2462, N2463);
nor NOR2_789 (N2539, N2467_t0, N2464_t0);
nor NOR2_790 (N2543, N2407_t1, N2470_t0);
nor NOR2_791 (N2544, N2470_t1, N2404_t1);
nor NOR2_792 (N2545, N2474, N2475);
nor NOR2_793 (N2548, N2476, N2477);
nor NOR2_794 (N2549, N2481, N2482);
nor NOR2_795 (N2552, N2486, N2487);
nor NOR2_796 (N2555, N2491, N2492);
nor NOR2_797 (N2558, N2496, N2497);
nor NOR2_798 (N2561, N2501, N2502);
nor NOR2_799 (N2564, N2506, N2507);
nor NOR2_800 (N2567, N2511, N2512);
nor NOR2_801 (N2570, N2516, N2517);
nor NOR2_802 (N2573, N2521, N2522);
nor NOR2_803 (N2576, N2526, N2527);
nor NOR2_804 (N2579, N2531, N2532);
nor NOR2_805 (N2582, N2536_t0, N2533_t0);
nor NOR2_806 (N2586, N2467_t1, N2539_t0);
nor NOR2_807 (N2587, N2539_t1, N2464_t1);
nor NOR2_808 (N2588, N2543, N2544);
nor NOR2_809 (N2591, N2545_t0, N1230_t0);
nor NOR2_810 (N2595, N2549_t0, N2478_t0);
nor NOR2_811 (N2599, N2552_t0, N2483_t0);
nor NOR2_812 (N2603, N2555_t0, N2488_t0);
nor NOR2_813 (N2607, N2558_t0, N2493_t0);
nor NOR2_814 (N2611, N2561_t0, N2498_t0);
nor NOR2_815 (N2615, N2564_t0, N2503_t0);
nor NOR2_816 (N2619, N2567_t0, N2508_t0);
nor NOR2_817 (N2623, N2570_t0, N2513_t0);
nor NOR2_818 (N2627, N2573_t0, N2518_t0);
nor NOR2_819 (N2631, N2576_t0, N2523_t0);
nor NOR2_820 (N2635, N2579_t0, N2528_t0);
nor NOR2_821 (N2639, N2536_t1, N2582_t0);
nor NOR2_822 (N2640, N2582_t1, N2533_t1);
nor NOR2_823 (N2641, N2586, N2587);
nor NOR2_824 (N2644, N2588_t0, N1182_t0);
nor NOR2_825 (N2648, N2545_t1, N2591_t0);
nor NOR2_826 (N2649, N2591_t1, N1230_t1);
nor NOR2_827 (N2650, N2410_t2, N2591_t2);
nor NOR2_828 (N2653, N2549_t1, N2595_t0);
nor NOR2_829 (N2654, N2595_t1, N2478_t1);
nor NOR2_830 (N2655, N2552_t1, N2599_t0);
nor NOR2_831 (N2656, N2599_t1, N2483_t1);
nor NOR2_832 (N2657, N2555_t1, N2603_t0);
nor NOR2_833 (N2658, N2603_t1, N2488_t1);
nor NOR2_834 (N2659, N2558_t1, N2607_t0);
nor NOR2_835 (N2660, N2607_t1, N2493_t1);
nor NOR2_836 (N2661, N2561_t1, N2611_t0);
nor NOR2_837 (N2662, N2611_t1, N2498_t1);
nor NOR2_838 (N2663, N2564_t1, N2615_t0);
nor NOR2_839 (N2664, N2615_t1, N2503_t1);
nor NOR2_840 (N2665, N2567_t1, N2619_t0);
nor NOR2_841 (N2666, N2619_t1, N2508_t1);
nor NOR2_842 (N2667, N2570_t1, N2623_t0);
nor NOR2_843 (N2668, N2623_t1, N2513_t1);
nor NOR2_844 (N2669, N2573_t1, N2627_t0);
nor NOR2_845 (N2670, N2627_t1, N2518_t1);
nor NOR2_846 (N2671, N2576_t1, N2631_t0);
nor NOR2_847 (N2672, N2631_t1, N2523_t1);
nor NOR2_848 (N2673, N2579_t1, N2635_t0);
nor NOR2_849 (N2674, N2635_t1, N2528_t1);
nor NOR2_850 (N2675, N2639, N2640);
nor NOR2_851 (N2678, N2641_t0, N1134_t0);
nor NOR2_852 (N2682, N2588_t1, N2644_t0);
nor NOR2_853 (N2683, N2644_t1, N1182_t1);
nor NOR2_854 (N2684, N2470_t2, N2644_t2);
nor NOR2_855 (N2687, N2648, N2649);
nor NOR2_856 (N2690, N1278_t0, N2650_t0);
nor NOR2_857 (N2694, N2653, N2654);
nor NOR2_858 (N2697, N2655, N2656);
nor NOR2_859 (N2700, N2657, N2658);
nor NOR2_860 (N2703, N2659, N2660);
nor NOR2_861 (N2706, N2661, N2662);
nor NOR2_862 (N2709, N2663, N2664);
nor NOR2_863 (N2712, N2665, N2666);
nor NOR2_864 (N2715, N2667, N2668);
nor NOR2_865 (N2718, N2669, N2670);
nor NOR2_866 (N2721, N2671, N2672);
nor NOR2_867 (N2724, N2673, N2674);
nor NOR2_868 (N2727, N2675_t0, N1086_t0);
nor NOR2_869 (N2731, N2641_t1, N2678_t0);
nor NOR2_870 (N2732, N2678_t1, N1134_t1);
nor NOR2_871 (N2733, N2539_t2, N2678_t2);
nor NOR2_872 (N2736, N2682, N2683);
nor NOR2_873 (N2739, N2687_t0, N2684_t0);
nor NOR2_874 (N2743, N1278_t1, N2690_t0);
nor NOR2_875 (N2744, N2690_t1, N2650_t1);
nor NOR2_876 (N2745, N2694_t0, N558_t0);
nor NOR2_877 (N2749, N2697_t0, N606_t0);
nor NOR2_878 (N2753, N2700_t0, N654_t0);
nor NOR2_879 (N2757, N2703_t0, N702_t0);
nor NOR2_880 (N2761, N2706_t0, N750_t0);
nor NOR2_881 (N2765, N2709_t0, N798_t0);
nor NOR2_882 (N2769, N2712_t0, N846_t0);
nor NOR2_883 (N2773, N2715_t0, N894_t0);
nor NOR2_884 (N2777, N2718_t0, N942_t0);
nor NOR2_885 (N2781, N2721_t0, N990_t0);
nor NOR2_886 (N2785, N2724_t0, N1038_t0);
nor NOR2_887 (N2789, N2675_t1, N2727_t0);
nor NOR2_888 (N2790, N2727_t1, N1086_t1);
nor NOR2_889 (N2791, N2582_t2, N2727_t2);
nor NOR2_890 (N2794, N2731, N2732);
nor NOR2_891 (N2797, N2736_t0, N2733_t0);
nor NOR2_892 (N2801, N2687_t1, N2739_t0);
nor NOR2_893 (N2802, N2739_t1, N2684_t1);
nor NOR2_894 (N2803, N2743, N2744);
nor NOR2_895 (N2806, N2694_t1, N2745_t0);
nor NOR2_896 (N2807, N2745_t1, N558_t1);
nor NOR2_897 (N2808, N2595_t2, N2745_t2);
nor NOR2_898 (N2811, N2697_t1, N2749_t0);
nor NOR2_899 (N2812, N2749_t1, N606_t1);
nor NOR2_900 (N2813, N2599_t2, N2749_t2);
nor NOR2_901 (N2816, N2700_t1, N2753_t0);
nor NOR2_902 (N2817, N2753_t1, N654_t1);
nor NOR2_903 (N2818, N2603_t2, N2753_t2);
nor NOR2_904 (N2821, N2703_t1, N2757_t0);
nor NOR2_905 (N2822, N2757_t1, N702_t1);
nor NOR2_906 (N2823, N2607_t2, N2757_t2);
nor NOR2_907 (N2826, N2706_t1, N2761_t0);
nor NOR2_908 (N2827, N2761_t1, N750_t1);
nor NOR2_909 (N2828, N2611_t2, N2761_t2);
nor NOR2_910 (N2831, N2709_t1, N2765_t0);
nor NOR2_911 (N2832, N2765_t1, N798_t1);
nor NOR2_912 (N2833, N2615_t2, N2765_t2);
nor NOR2_913 (N2836, N2712_t1, N2769_t0);
nor NOR2_914 (N2837, N2769_t1, N846_t1);
nor NOR2_915 (N2838, N2619_t2, N2769_t2);
nor NOR2_916 (N2841, N2715_t1, N2773_t0);
nor NOR2_917 (N2842, N2773_t1, N894_t1);
nor NOR2_918 (N2843, N2623_t2, N2773_t2);
nor NOR2_919 (N2846, N2718_t1, N2777_t0);
nor NOR2_920 (N2847, N2777_t1, N942_t1);
nor NOR2_921 (N2848, N2627_t2, N2777_t2);
nor NOR2_922 (N2851, N2721_t1, N2781_t0);
nor NOR2_923 (N2852, N2781_t1, N990_t1);
nor NOR2_924 (N2853, N2631_t2, N2781_t2);
nor NOR2_925 (N2856, N2724_t1, N2785_t0);
nor NOR2_926 (N2857, N2785_t1, N1038_t1);
nor NOR2_927 (N2858, N2635_t2, N2785_t2);
nor NOR2_928 (N2861, N2789, N2790);
nor NOR2_929 (N2864, N2794_t0, N2791_t0);
nor NOR2_930 (N2868, N2736_t1, N2797_t0);
nor NOR2_931 (N2869, N2797_t1, N2733_t1);
nor NOR2_932 (N2870, N2801, N2802);
nor NOR2_933 (N2873, N2803_t0, N1233_t0);
nor NOR2_934 (N2877, N2806, N2807);
nor NOR2_935 (N2878, N2811, N2812);
nor NOR2_936 (N2881, N2816, N2817);
nor NOR2_937 (N2884, N2821, N2822);
nor NOR2_938 (N2887, N2826, N2827);
nor NOR2_939 (N2890, N2831, N2832);
nor NOR2_940 (N2893, N2836, N2837);
nor NOR2_941 (N2896, N2841, N2842);
nor NOR2_942 (N2899, N2846, N2847);
nor NOR2_943 (N2902, N2851, N2852);
nor NOR2_944 (N2905, N2856, N2857);
nor NOR2_945 (N2908, N2861_t0, N2858_t0);
nor NOR2_946 (N2912, N2794_t1, N2864_t0);
nor NOR2_947 (N2913, N2864_t1, N2791_t1);
nor NOR2_948 (N2914, N2868, N2869);
nor NOR2_949 (N2917, N2870_t0, N1185_t0);
nor NOR2_950 (N2921, N2803_t1, N2873_t0);
nor NOR2_951 (N2922, N2873_t1, N1233_t1);
nor NOR2_952 (N2923, N2690_t2, N2873_t2);
nor NOR2_953 (N2926, N2878_t0, N2808_t0);
nor NOR2_954 (N2930, N2881_t0, N2813_t0);
nor NOR2_955 (N2934, N2884_t0, N2818_t0);
nor NOR2_956 (N2938, N2887_t0, N2823_t0);
nor NOR2_957 (N2942, N2890_t0, N2828_t0);
nor NOR2_958 (N2946, N2893_t0, N2833_t0);
nor NOR2_959 (N2950, N2896_t0, N2838_t0);
nor NOR2_960 (N2954, N2899_t0, N2843_t0);
nor NOR2_961 (N2958, N2902_t0, N2848_t0);
nor NOR2_962 (N2962, N2905_t0, N2853_t0);
nor NOR2_963 (N2966, N2861_t1, N2908_t0);
nor NOR2_964 (N2967, N2908_t1, N2858_t1);
nor NOR2_965 (N2968, N2912, N2913);
nor NOR2_966 (N2971, N2914_t0, N1137_t0);
nor NOR2_967 (N2975, N2870_t1, N2917_t0);
nor NOR2_968 (N2976, N2917_t1, N1185_t1);
nor NOR2_969 (N2977, N2739_t2, N2917_t2);
nor NOR2_970 (N2980, N2921, N2922);
nor NOR2_971 (N2983, N1281_t0, N2923_t0);
nor NOR2_972 (N2987, N2878_t1, N2926_t0);
nor NOR2_973 (N2988, N2926_t1, N2808_t1);
nor NOR2_974 (N2989, N2881_t1, N2930_t0);
nor NOR2_975 (N2990, N2930_t1, N2813_t1);
nor NOR2_976 (N2991, N2884_t1, N2934_t0);
nor NOR2_977 (N2992, N2934_t1, N2818_t1);
nor NOR2_978 (N2993, N2887_t1, N2938_t0);
nor NOR2_979 (N2994, N2938_t1, N2823_t1);
nor NOR2_980 (N2995, N2890_t1, N2942_t0);
nor NOR2_981 (N2996, N2942_t1, N2828_t1);
nor NOR2_982 (N2997, N2893_t1, N2946_t0);
nor NOR2_983 (N2998, N2946_t1, N2833_t1);
nor NOR2_984 (N2999, N2896_t1, N2950_t0);
nor NOR2_985 (N3000, N2950_t1, N2838_t1);
nor NOR2_986 (N3001, N2899_t1, N2954_t0);
nor NOR2_987 (N3002, N2954_t1, N2843_t1);
nor NOR2_988 (N3003, N2902_t1, N2958_t0);
nor NOR2_989 (N3004, N2958_t1, N2848_t1);
nor NOR2_990 (N3005, N2905_t1, N2962_t0);
nor NOR2_991 (N3006, N2962_t1, N2853_t1);
nor NOR2_992 (N3007, N2966, N2967);
nor NOR2_993 (N3010, N2968_t0, N1089_t0);
nor NOR2_994 (N3014, N2914_t1, N2971_t0);
nor NOR2_995 (N3015, N2971_t1, N1137_t1);
nor NOR2_996 (N3016, N2797_t2, N2971_t2);
nor NOR2_997 (N3019, N2975, N2976);
nor NOR2_998 (N3022, N2980_t0, N2977_t0);
nor NOR2_999 (N3026, N1281_t1, N2983_t0);
nor NOR2_1000 (N3027, N2983_t1, N2923_t1);
nor NOR2_1001 (N3028, N2987, N2988);
nor NOR2_1002 (N3031, N2989, N2990);
nor NOR2_1003 (N3034, N2991, N2992);
nor NOR2_1004 (N3037, N2993, N2994);
nor NOR2_1005 (N3040, N2995, N2996);
nor NOR2_1006 (N3043, N2997, N2998);
nor NOR2_1007 (N3046, N2999, N3000);
nor NOR2_1008 (N3049, N3001, N3002);
nor NOR2_1009 (N3052, N3003, N3004);
nor NOR2_1010 (N3055, N3005, N3006);
nor NOR2_1011 (N3058, N3007_t0, N1041_t0);
nor NOR2_1012 (N3062, N2968_t1, N3010_t0);
nor NOR2_1013 (N3063, N3010_t1, N1089_t1);
nor NOR2_1014 (N3064, N2864_t2, N3010_t2);
nor NOR2_1015 (N3067, N3014, N3015);
nor NOR2_1016 (N3070, N3019_t0, N3016_t0);
nor NOR2_1017 (N3074, N2980_t1, N3022_t0);
nor NOR2_1018 (N3075, N3022_t1, N2977_t1);
nor NOR2_1019 (N3076, N3026, N3027);
nor NOR2_1020 (N3079, N3028_t0, N561_t0);
nor NOR2_1021 (N3083, N3031_t0, N609_t0);
nor NOR2_1022 (N3087, N3034_t0, N657_t0);
nor NOR2_1023 (N3091, N3037_t0, N705_t0);
nor NOR2_1024 (N3095, N3040_t0, N753_t0);
nor NOR2_1025 (N3099, N3043_t0, N801_t0);
nor NOR2_1026 (N3103, N3046_t0, N849_t0);
nor NOR2_1027 (N3107, N3049_t0, N897_t0);
nor NOR2_1028 (N3111, N3052_t0, N945_t0);
nor NOR2_1029 (N3115, N3055_t0, N993_t0);
nor NOR2_1030 (N3119, N3007_t1, N3058_t0);
nor NOR2_1031 (N3120, N3058_t1, N1041_t1);
nor NOR2_1032 (N3121, N2908_t2, N3058_t2);
nor NOR2_1033 (N3124, N3062, N3063);
nor NOR2_1034 (N3127, N3067_t0, N3064_t0);
nor NOR2_1035 (N3131, N3019_t1, N3070_t0);
nor NOR2_1036 (N3132, N3070_t1, N3016_t1);
nor NOR2_1037 (N3133, N3074, N3075);
nor NOR2_1038 (N3136, N3076_t0, N1236_t0);
nor NOR2_1039 (N3140, N3028_t1, N3079_t0);
nor NOR2_1040 (N3141, N3079_t1, N561_t1);
nor NOR2_1041 (N3142, N2926_t2, N3079_t2);
nor NOR2_1042 (N3145, N3031_t1, N3083_t0);
nor NOR2_1043 (N3146, N3083_t1, N609_t1);
nor NOR2_1044 (N3147, N2930_t2, N3083_t2);
nor NOR2_1045 (N3150, N3034_t1, N3087_t0);
nor NOR2_1046 (N3151, N3087_t1, N657_t1);
nor NOR2_1047 (N3152, N2934_t2, N3087_t2);
nor NOR2_1048 (N3155, N3037_t1, N3091_t0);
nor NOR2_1049 (N3156, N3091_t1, N705_t1);
nor NOR2_1050 (N3157, N2938_t2, N3091_t2);
nor NOR2_1051 (N3160, N3040_t1, N3095_t0);
nor NOR2_1052 (N3161, N3095_t1, N753_t1);
nor NOR2_1053 (N3162, N2942_t2, N3095_t2);
nor NOR2_1054 (N3165, N3043_t1, N3099_t0);
nor NOR2_1055 (N3166, N3099_t1, N801_t1);
nor NOR2_1056 (N3167, N2946_t2, N3099_t2);
nor NOR2_1057 (N3170, N3046_t1, N3103_t0);
nor NOR2_1058 (N3171, N3103_t1, N849_t1);
nor NOR2_1059 (N3172, N2950_t2, N3103_t2);
nor NOR2_1060 (N3175, N3049_t1, N3107_t0);
nor NOR2_1061 (N3176, N3107_t1, N897_t1);
nor NOR2_1062 (N3177, N2954_t2, N3107_t2);
nor NOR2_1063 (N3180, N3052_t1, N3111_t0);
nor NOR2_1064 (N3181, N3111_t1, N945_t1);
nor NOR2_1065 (N3182, N2958_t2, N3111_t2);
nor NOR2_1066 (N3185, N3055_t1, N3115_t0);
nor NOR2_1067 (N3186, N3115_t1, N993_t1);
nor NOR2_1068 (N3187, N2962_t2, N3115_t2);
nor NOR2_1069 (N3190, N3119, N3120);
nor NOR2_1070 (N3193, N3124_t0, N3121_t0);
nor NOR2_1071 (N3197, N3067_t1, N3127_t0);
nor NOR2_1072 (N3198, N3127_t1, N3064_t1);
nor NOR2_1073 (N3199, N3131, N3132);
nor NOR2_1074 (N3202, N3133_t0, N1188_t0);
nor NOR2_1075 (N3206, N3076_t1, N3136_t0);
nor NOR2_1076 (N3207, N3136_t1, N1236_t1);
nor NOR2_1077 (N3208, N2983_t2, N3136_t2);
nor NOR2_1078 (N3211, N3140, N3141);
nor NOR2_1079 (N3212, N3145, N3146);
nor NOR2_1080 (N3215, N3150, N3151);
nor NOR2_1081 (N3218, N3155, N3156);
nor NOR2_1082 (N3221, N3160, N3161);
nor NOR2_1083 (N3224, N3165, N3166);
nor NOR2_1084 (N3227, N3170, N3171);
nor NOR2_1085 (N3230, N3175, N3176);
nor NOR2_1086 (N3233, N3180, N3181);
nor NOR2_1087 (N3236, N3185, N3186);
nor NOR2_1088 (N3239, N3190_t0, N3187_t0);
nor NOR2_1089 (N3243, N3124_t1, N3193_t0);
nor NOR2_1090 (N3244, N3193_t1, N3121_t1);
nor NOR2_1091 (N3245, N3197, N3198);
nor NOR2_1092 (N3248, N3199_t0, N1140_t0);
nor NOR2_1093 (N3252, N3133_t1, N3202_t0);
nor NOR2_1094 (N3253, N3202_t1, N1188_t1);
nor NOR2_1095 (N3254, N3022_t2, N3202_t2);
nor NOR2_1096 (N3257, N3206, N3207);
nor NOR2_1097 (N3260, N1284_t0, N3208_t0);
nor NOR2_1098 (N3264, N3212_t0, N3142_t0);
nor NOR2_1099 (N3268, N3215_t0, N3147_t0);
nor NOR2_1100 (N3272, N3218_t0, N3152_t0);
nor NOR2_1101 (N3276, N3221_t0, N3157_t0);
nor NOR2_1102 (N3280, N3224_t0, N3162_t0);
nor NOR2_1103 (N3284, N3227_t0, N3167_t0);
nor NOR2_1104 (N3288, N3230_t0, N3172_t0);
nor NOR2_1105 (N3292, N3233_t0, N3177_t0);
nor NOR2_1106 (N3296, N3236_t0, N3182_t0);
nor NOR2_1107 (N3300, N3190_t1, N3239_t0);
nor NOR2_1108 (N3301, N3239_t1, N3187_t1);
nor NOR2_1109 (N3302, N3243, N3244);
nor NOR2_1110 (N3305, N3245_t0, N1092_t0);
nor NOR2_1111 (N3309, N3199_t1, N3248_t0);
nor NOR2_1112 (N3310, N3248_t1, N1140_t1);
nor NOR2_1113 (N3311, N3070_t2, N3248_t2);
nor NOR2_1114 (N3314, N3252, N3253);
nor NOR2_1115 (N3317, N3257_t0, N3254_t0);
nor NOR2_1116 (N3321, N1284_t1, N3260_t0);
nor NOR2_1117 (N3322, N3260_t1, N3208_t1);
nor NOR2_1118 (N3323, N3212_t1, N3264_t0);
nor NOR2_1119 (N3324, N3264_t1, N3142_t1);
nor NOR2_1120 (N3325, N3215_t1, N3268_t0);
nor NOR2_1121 (N3326, N3268_t1, N3147_t1);
nor NOR2_1122 (N3327, N3218_t1, N3272_t0);
nor NOR2_1123 (N3328, N3272_t1, N3152_t1);
nor NOR2_1124 (N3329, N3221_t1, N3276_t0);
nor NOR2_1125 (N3330, N3276_t1, N3157_t1);
nor NOR2_1126 (N3331, N3224_t1, N3280_t0);
nor NOR2_1127 (N3332, N3280_t1, N3162_t1);
nor NOR2_1128 (N3333, N3227_t1, N3284_t0);
nor NOR2_1129 (N3334, N3284_t1, N3167_t1);
nor NOR2_1130 (N3335, N3230_t1, N3288_t0);
nor NOR2_1131 (N3336, N3288_t1, N3172_t1);
nor NOR2_1132 (N3337, N3233_t1, N3292_t0);
nor NOR2_1133 (N3338, N3292_t1, N3177_t1);
nor NOR2_1134 (N3339, N3236_t1, N3296_t0);
nor NOR2_1135 (N3340, N3296_t1, N3182_t1);
nor NOR2_1136 (N3341, N3300, N3301);
nor NOR2_1137 (N3344, N3302_t0, N1044_t0);
nor NOR2_1138 (N3348, N3245_t1, N3305_t0);
nor NOR2_1139 (N3349, N3305_t1, N1092_t1);
nor NOR2_1140 (N3350, N3127_t2, N3305_t2);
nor NOR2_1141 (N3353, N3309, N3310);
nor NOR2_1142 (N3356, N3314_t0, N3311_t0);
nor NOR2_1143 (N3360, N3257_t1, N3317_t0);
nor NOR2_1144 (N3361, N3317_t1, N3254_t1);
nor NOR2_1145 (N3362, N3321, N3322);
nor NOR2_1146 (N3365, N3323, N3324);
nor NOR2_1147 (N3368, N3325, N3326);
nor NOR2_1148 (N3371, N3327, N3328);
nor NOR2_1149 (N3374, N3329, N3330);
nor NOR2_1150 (N3377, N3331, N3332);
nor NOR2_1151 (N3380, N3333, N3334);
nor NOR2_1152 (N3383, N3335, N3336);
nor NOR2_1153 (N3386, N3337, N3338);
nor NOR2_1154 (N3389, N3339, N3340);
nor NOR2_1155 (N3392, N3341_t0, N996_t0);
nor NOR2_1156 (N3396, N3302_t1, N3344_t0);
nor NOR2_1157 (N3397, N3344_t1, N1044_t1);
nor NOR2_1158 (N3398, N3193_t2, N3344_t2);
nor NOR2_1159 (N3401, N3348, N3349);
nor NOR2_1160 (N3404, N3353_t0, N3350_t0);
nor NOR2_1161 (N3408, N3314_t1, N3356_t0);
nor NOR2_1162 (N3409, N3356_t1, N3311_t1);
nor NOR2_1163 (N3410, N3360, N3361);
nor NOR2_1164 (N3413, N3362_t0, N1239_t0);
nor NOR2_1165 (N3417, N3365_t0, N564_t0);
nor NOR2_1166 (N3421, N3368_t0, N612_t0);
nor NOR2_1167 (N3425, N3371_t0, N660_t0);
nor NOR2_1168 (N3429, N3374_t0, N708_t0);
nor NOR2_1169 (N3433, N3377_t0, N756_t0);
nor NOR2_1170 (N3437, N3380_t0, N804_t0);
nor NOR2_1171 (N3441, N3383_t0, N852_t0);
nor NOR2_1172 (N3445, N3386_t0, N900_t0);
nor NOR2_1173 (N3449, N3389_t0, N948_t0);
nor NOR2_1174 (N3453, N3341_t1, N3392_t0);
nor NOR2_1175 (N3454, N3392_t1, N996_t1);
nor NOR2_1176 (N3455, N3239_t2, N3392_t2);
nor NOR2_1177 (N3458, N3396, N3397);
nor NOR2_1178 (N3461, N3401_t0, N3398_t0);
nor NOR2_1179 (N3465, N3353_t1, N3404_t0);
nor NOR2_1180 (N3466, N3404_t1, N3350_t1);
nor NOR2_1181 (N3467, N3408, N3409);
nor NOR2_1182 (N3470, N3410_t0, N1191_t0);
nor NOR2_1183 (N3474, N3362_t1, N3413_t0);
nor NOR2_1184 (N3475, N3413_t1, N1239_t1);
nor NOR2_1185 (N3476, N3260_t2, N3413_t2);
nor NOR2_1186 (N3479, N3365_t1, N3417_t0);
nor NOR2_1187 (N3480, N3417_t1, N564_t1);
nor NOR2_1188 (N3481, N3264_t2, N3417_t2);
nor NOR2_1189 (N3484, N3368_t1, N3421_t0);
nor NOR2_1190 (N3485, N3421_t1, N612_t1);
nor NOR2_1191 (N3486, N3268_t2, N3421_t2);
nor NOR2_1192 (N3489, N3371_t1, N3425_t0);
nor NOR2_1193 (N3490, N3425_t1, N660_t1);
nor NOR2_1194 (N3491, N3272_t2, N3425_t2);
nor NOR2_1195 (N3494, N3374_t1, N3429_t0);
nor NOR2_1196 (N3495, N3429_t1, N708_t1);
nor NOR2_1197 (N3496, N3276_t2, N3429_t2);
nor NOR2_1198 (N3499, N3377_t1, N3433_t0);
nor NOR2_1199 (N3500, N3433_t1, N756_t1);
nor NOR2_1200 (N3501, N3280_t2, N3433_t2);
nor NOR2_1201 (N3504, N3380_t1, N3437_t0);
nor NOR2_1202 (N3505, N3437_t1, N804_t1);
nor NOR2_1203 (N3506, N3284_t2, N3437_t2);
nor NOR2_1204 (N3509, N3383_t1, N3441_t0);
nor NOR2_1205 (N3510, N3441_t1, N852_t1);
nor NOR2_1206 (N3511, N3288_t2, N3441_t2);
nor NOR2_1207 (N3514, N3386_t1, N3445_t0);
nor NOR2_1208 (N3515, N3445_t1, N900_t1);
nor NOR2_1209 (N3516, N3292_t2, N3445_t2);
nor NOR2_1210 (N3519, N3389_t1, N3449_t0);
nor NOR2_1211 (N3520, N3449_t1, N948_t1);
nor NOR2_1212 (N3521, N3296_t2, N3449_t2);
nor NOR2_1213 (N3524, N3453, N3454);
nor NOR2_1214 (N3527, N3458_t0, N3455_t0);
nor NOR2_1215 (N3531, N3401_t1, N3461_t0);
nor NOR2_1216 (N3532, N3461_t1, N3398_t1);
nor NOR2_1217 (N3533, N3465, N3466);
nor NOR2_1218 (N3536, N3467_t0, N1143_t0);
nor NOR2_1219 (N3540, N3410_t1, N3470_t0);
nor NOR2_1220 (N3541, N3470_t1, N1191_t1);
nor NOR2_1221 (N3542, N3317_t2, N3470_t2);
nor NOR2_1222 (N3545, N3474, N3475);
nor NOR2_1223 (N3548, N1287_t0, N3476_t0);
nor NOR2_1224 (N3552, N3479, N3480);
nor NOR2_1225 (N3553, N3484, N3485);
nor NOR2_1226 (N3556, N3489, N3490);
nor NOR2_1227 (N3559, N3494, N3495);
nor NOR2_1228 (N3562, N3499, N3500);
nor NOR2_1229 (N3565, N3504, N3505);
nor NOR2_1230 (N3568, N3509, N3510);
nor NOR2_1231 (N3571, N3514, N3515);
nor NOR2_1232 (N3574, N3519, N3520);
nor NOR2_1233 (N3577, N3524_t0, N3521_t0);
nor NOR2_1234 (N3581, N3458_t1, N3527_t0);
nor NOR2_1235 (N3582, N3527_t1, N3455_t1);
nor NOR2_1236 (N3583, N3531, N3532);
nor NOR2_1237 (N3586, N3533_t0, N1095_t0);
nor NOR2_1238 (N3590, N3467_t1, N3536_t0);
nor NOR2_1239 (N3591, N3536_t1, N1143_t1);
nor NOR2_1240 (N3592, N3356_t2, N3536_t2);
nor NOR2_1241 (N3595, N3540, N3541);
nor NOR2_1242 (N3598, N3545_t0, N3542_t0);
nor NOR2_1243 (N3602, N1287_t1, N3548_t0);
nor NOR2_1244 (N3603, N3548_t1, N3476_t1);
nor NOR2_1245 (N3604, N3553_t0, N3481_t0);
nor NOR2_1246 (N3608, N3556_t0, N3486_t0);
nor NOR2_1247 (N3612, N3559_t0, N3491_t0);
nor NOR2_1248 (N3616, N3562_t0, N3496_t0);
nor NOR2_1249 (N3620, N3565_t0, N3501_t0);
nor NOR2_1250 (N3624, N3568_t0, N3506_t0);
nor NOR2_1251 (N3628, N3571_t0, N3511_t0);
nor NOR2_1252 (N3632, N3574_t0, N3516_t0);
nor NOR2_1253 (N3636, N3524_t1, N3577_t0);
nor NOR2_1254 (N3637, N3577_t1, N3521_t1);
nor NOR2_1255 (N3638, N3581, N3582);
nor NOR2_1256 (N3641, N3583_t0, N1047_t0);
nor NOR2_1257 (N3645, N3533_t1, N3586_t0);
nor NOR2_1258 (N3646, N3586_t1, N1095_t1);
nor NOR2_1259 (N3647, N3404_t2, N3586_t2);
nor NOR2_1260 (N3650, N3590, N3591);
nor NOR2_1261 (N3653, N3595_t0, N3592_t0);
nor NOR2_1262 (N3657, N3545_t1, N3598_t0);
nor NOR2_1263 (N3658, N3598_t1, N3542_t1);
nor NOR2_1264 (N3659, N3602, N3603);
nor NOR2_1265 (N3662, N3553_t1, N3604_t0);
nor NOR2_1266 (N3663, N3604_t1, N3481_t1);
nor NOR2_1267 (N3664, N3556_t1, N3608_t0);
nor NOR2_1268 (N3665, N3608_t1, N3486_t1);
nor NOR2_1269 (N3666, N3559_t1, N3612_t0);
nor NOR2_1270 (N3667, N3612_t1, N3491_t1);
nor NOR2_1271 (N3668, N3562_t1, N3616_t0);
nor NOR2_1272 (N3669, N3616_t1, N3496_t1);
nor NOR2_1273 (N3670, N3565_t1, N3620_t0);
nor NOR2_1274 (N3671, N3620_t1, N3501_t1);
nor NOR2_1275 (N3672, N3568_t1, N3624_t0);
nor NOR2_1276 (N3673, N3624_t1, N3506_t1);
nor NOR2_1277 (N3674, N3571_t1, N3628_t0);
nor NOR2_1278 (N3675, N3628_t1, N3511_t1);
nor NOR2_1279 (N3676, N3574_t1, N3632_t0);
nor NOR2_1280 (N3677, N3632_t1, N3516_t1);
nor NOR2_1281 (N3678, N3636, N3637);
nor NOR2_1282 (N3681, N3638_t0, N999_t0);
nor NOR2_1283 (N3685, N3583_t1, N3641_t0);
nor NOR2_1284 (N3686, N3641_t1, N1047_t1);
nor NOR2_1285 (N3687, N3461_t2, N3641_t2);
nor NOR2_1286 (N3690, N3645, N3646);
nor NOR2_1287 (N3693, N3650_t0, N3647_t0);
nor NOR2_1288 (N3697, N3595_t1, N3653_t0);
nor NOR2_1289 (N3698, N3653_t1, N3592_t1);
nor NOR2_1290 (N3699, N3657, N3658);
nor NOR2_1291 (N3702, N3659_t0, N1242_t0);
nor NOR2_1292 (N3706, N3662, N3663);
nor NOR2_1293 (N3709, N3664, N3665);
nor NOR2_1294 (N3712, N3666, N3667);
nor NOR2_1295 (N3715, N3668, N3669);
nor NOR2_1296 (N3718, N3670, N3671);
nor NOR2_1297 (N3721, N3672, N3673);
nor NOR2_1298 (N3724, N3674, N3675);
nor NOR2_1299 (N3727, N3676, N3677);
nor NOR2_1300 (N3730, N3678_t0, N951_t0);
nor NOR2_1301 (N3734, N3638_t1, N3681_t0);
nor NOR2_1302 (N3735, N3681_t1, N999_t1);
nor NOR2_1303 (N3736, N3527_t2, N3681_t2);
nor NOR2_1304 (N3739, N3685, N3686);
nor NOR2_1305 (N3742, N3690_t0, N3687_t0);
nor NOR2_1306 (N3746, N3650_t1, N3693_t0);
nor NOR2_1307 (N3747, N3693_t1, N3647_t1);
nor NOR2_1308 (N3748, N3697, N3698);
nor NOR2_1309 (N3751, N3699_t0, N1194_t0);
nor NOR2_1310 (N3755, N3659_t1, N3702_t0);
nor NOR2_1311 (N3756, N3702_t1, N1242_t1);
nor NOR2_1312 (N3757, N3548_t2, N3702_t2);
nor NOR2_1313 (N3760, N3706_t0, N567_t0);
nor NOR2_1314 (N3764, N3709_t0, N615_t0);
nor NOR2_1315 (N3768, N3712_t0, N663_t0);
nor NOR2_1316 (N3772, N3715_t0, N711_t0);
nor NOR2_1317 (N3776, N3718_t0, N759_t0);
nor NOR2_1318 (N3780, N3721_t0, N807_t0);
nor NOR2_1319 (N3784, N3724_t0, N855_t0);
nor NOR2_1320 (N3788, N3727_t0, N903_t0);
nor NOR2_1321 (N3792, N3678_t1, N3730_t0);
nor NOR2_1322 (N3793, N3730_t1, N951_t1);
nor NOR2_1323 (N3794, N3577_t2, N3730_t2);
nor NOR2_1324 (N3797, N3734, N3735);
nor NOR2_1325 (N3800, N3739_t0, N3736_t0);
nor NOR2_1326 (N3804, N3690_t1, N3742_t0);
nor NOR2_1327 (N3805, N3742_t1, N3687_t1);
nor NOR2_1328 (N3806, N3746, N3747);
nor NOR2_1329 (N3809, N3748_t0, N1146_t0);
nor NOR2_1330 (N3813, N3699_t1, N3751_t0);
nor NOR2_1331 (N3814, N3751_t1, N1194_t1);
nor NOR2_1332 (N3815, N3598_t2, N3751_t2);
nor NOR2_1333 (N3818, N3755, N3756);
nor NOR2_1334 (N3821, N1290_t0, N3757_t0);
nor NOR2_1335 (N3825, N3706_t1, N3760_t0);
nor NOR2_1336 (N3826, N3760_t1, N567_t1);
nor NOR2_1337 (N3827, N3604_t2, N3760_t2);
nor NOR2_1338 (N3830, N3709_t1, N3764_t0);
nor NOR2_1339 (N3831, N3764_t1, N615_t1);
nor NOR2_1340 (N3832, N3608_t2, N3764_t2);
nor NOR2_1341 (N3835, N3712_t1, N3768_t0);
nor NOR2_1342 (N3836, N3768_t1, N663_t1);
nor NOR2_1343 (N3837, N3612_t2, N3768_t2);
nor NOR2_1344 (N3840, N3715_t1, N3772_t0);
nor NOR2_1345 (N3841, N3772_t1, N711_t1);
nor NOR2_1346 (N3842, N3616_t2, N3772_t2);
nor NOR2_1347 (N3845, N3718_t1, N3776_t0);
nor NOR2_1348 (N3846, N3776_t1, N759_t1);
nor NOR2_1349 (N3847, N3620_t2, N3776_t2);
nor NOR2_1350 (N3850, N3721_t1, N3780_t0);
nor NOR2_1351 (N3851, N3780_t1, N807_t1);
nor NOR2_1352 (N3852, N3624_t2, N3780_t2);
nor NOR2_1353 (N3855, N3724_t1, N3784_t0);
nor NOR2_1354 (N3856, N3784_t1, N855_t1);
nor NOR2_1355 (N3857, N3628_t2, N3784_t2);
nor NOR2_1356 (N3860, N3727_t1, N3788_t0);
nor NOR2_1357 (N3861, N3788_t1, N903_t1);
nor NOR2_1358 (N3862, N3632_t2, N3788_t2);
nor NOR2_1359 (N3865, N3792, N3793);
nor NOR2_1360 (N3868, N3797_t0, N3794_t0);
nor NOR2_1361 (N3872, N3739_t1, N3800_t0);
nor NOR2_1362 (N3873, N3800_t1, N3736_t1);
nor NOR2_1363 (N3874, N3804, N3805);
nor NOR2_1364 (N3877, N3806_t0, N1098_t0);
nor NOR2_1365 (N3881, N3748_t1, N3809_t0);
nor NOR2_1366 (N3882, N3809_t1, N1146_t1);
nor NOR2_1367 (N3883, N3653_t2, N3809_t2);
nor NOR2_1368 (N3886, N3813, N3814);
nor NOR2_1369 (N3889, N3818_t0, N3815_t0);
nor NOR2_1370 (N3893, N1290_t1, N3821_t0);
nor NOR2_1371 (N3894, N3821_t1, N3757_t1);
nor NOR2_1372 (N3895, N3825, N3826);
nor NOR2_1373 (N3896, N3830, N3831);
nor NOR2_1374 (N3899, N3835, N3836);
nor NOR2_1375 (N3902, N3840, N3841);
nor NOR2_1376 (N3905, N3845, N3846);
nor NOR2_1377 (N3908, N3850, N3851);
nor NOR2_1378 (N3911, N3855, N3856);
nor NOR2_1379 (N3914, N3860, N3861);
nor NOR2_1380 (N3917, N3865_t0, N3862_t0);
nor NOR2_1381 (N3921, N3797_t1, N3868_t0);
nor NOR2_1382 (N3922, N3868_t1, N3794_t1);
nor NOR2_1383 (N3923, N3872, N3873);
nor NOR2_1384 (N3926, N3874_t0, N1050_t0);
nor NOR2_1385 (N3930, N3806_t1, N3877_t0);
nor NOR2_1386 (N3931, N3877_t1, N1098_t1);
nor NOR2_1387 (N3932, N3693_t2, N3877_t2);
nor NOR2_1388 (N3935, N3881, N3882);
nor NOR2_1389 (N3938, N3886_t0, N3883_t0);
nor NOR2_1390 (N3942, N3818_t1, N3889_t0);
nor NOR2_1391 (N3943, N3889_t1, N3815_t1);
nor NOR2_1392 (N3944, N3893, N3894);
nor NOR2_1393 (N3947, N3896_t0, N3827_t0);
nor NOR2_1394 (N3951, N3899_t0, N3832_t0);
nor NOR2_1395 (N3955, N3902_t0, N3837_t0);
nor NOR2_1396 (N3959, N3905_t0, N3842_t0);
nor NOR2_1397 (N3963, N3908_t0, N3847_t0);
nor NOR2_1398 (N3967, N3911_t0, N3852_t0);
nor NOR2_1399 (N3971, N3914_t0, N3857_t0);
nor NOR2_1400 (N3975, N3865_t1, N3917_t0);
nor NOR2_1401 (N3976, N3917_t1, N3862_t1);
nor NOR2_1402 (N3977, N3921, N3922);
nor NOR2_1403 (N3980, N3923_t0, N1002_t0);
nor NOR2_1404 (N3984, N3874_t1, N3926_t0);
nor NOR2_1405 (N3985, N3926_t1, N1050_t1);
nor NOR2_1406 (N3986, N3742_t2, N3926_t2);
nor NOR2_1407 (N3989, N3930, N3931);
nor NOR2_1408 (N3992, N3935_t0, N3932_t0);
nor NOR2_1409 (N3996, N3886_t1, N3938_t0);
nor NOR2_1410 (N3997, N3938_t1, N3883_t1);
nor NOR2_1411 (N3998, N3942, N3943);
nor NOR2_1412 (N4001, N3944_t0, N1245_t0);
nor NOR2_1413 (N4005, N3896_t1, N3947_t0);
nor NOR2_1414 (N4006, N3947_t1, N3827_t1);
nor NOR2_1415 (N4007, N3899_t1, N3951_t0);
nor NOR2_1416 (N4008, N3951_t1, N3832_t1);
nor NOR2_1417 (N4009, N3902_t1, N3955_t0);
nor NOR2_1418 (N4010, N3955_t1, N3837_t1);
nor NOR2_1419 (N4011, N3905_t1, N3959_t0);
nor NOR2_1420 (N4012, N3959_t1, N3842_t1);
nor NOR2_1421 (N4013, N3908_t1, N3963_t0);
nor NOR2_1422 (N4014, N3963_t1, N3847_t1);
nor NOR2_1423 (N4015, N3911_t1, N3967_t0);
nor NOR2_1424 (N4016, N3967_t1, N3852_t1);
nor NOR2_1425 (N4017, N3914_t1, N3971_t0);
nor NOR2_1426 (N4018, N3971_t1, N3857_t1);
nor NOR2_1427 (N4019, N3975, N3976);
nor NOR2_1428 (N4022, N3977_t0, N954_t0);
nor NOR2_1429 (N4026, N3923_t1, N3980_t0);
nor NOR2_1430 (N4027, N3980_t1, N1002_t1);
nor NOR2_1431 (N4028, N3800_t2, N3980_t2);
nor NOR2_1432 (N4031, N3984, N3985);
nor NOR2_1433 (N4034, N3989_t0, N3986_t0);
nor NOR2_1434 (N4038, N3935_t1, N3992_t0);
nor NOR2_1435 (N4039, N3992_t1, N3932_t1);
nor NOR2_1436 (N4040, N3996, N3997);
nor NOR2_1437 (N4043, N3998_t0, N1197_t0);
nor NOR2_1438 (N4047, N3944_t1, N4001_t0);
nor NOR2_1439 (N4048, N4001_t1, N1245_t1);
nor NOR2_1440 (N4049, N3821_t2, N4001_t2);
nor NOR2_1441 (N4052, N4005, N4006);
nor NOR2_1442 (N4055, N4007, N4008);
nor NOR2_1443 (N4058, N4009, N4010);
nor NOR2_1444 (N4061, N4011, N4012);
nor NOR2_1445 (N4064, N4013, N4014);
nor NOR2_1446 (N4067, N4015, N4016);
nor NOR2_1447 (N4070, N4017, N4018);
nor NOR2_1448 (N4073, N4019_t0, N906_t0);
nor NOR2_1449 (N4077, N3977_t1, N4022_t0);
nor NOR2_1450 (N4078, N4022_t1, N954_t1);
nor NOR2_1451 (N4079, N3868_t2, N4022_t2);
nor NOR2_1452 (N4082, N4026, N4027);
nor NOR2_1453 (N4085, N4031_t0, N4028_t0);
nor NOR2_1454 (N4089, N3989_t1, N4034_t0);
nor NOR2_1455 (N4090, N4034_t1, N3986_t1);
nor NOR2_1456 (N4091, N4038, N4039);
nor NOR2_1457 (N4094, N4040_t0, N1149_t0);
nor NOR2_1458 (N4098, N3998_t1, N4043_t0);
nor NOR2_1459 (N4099, N4043_t1, N1197_t1);
nor NOR2_1460 (N4100, N3889_t2, N4043_t2);
nor NOR2_1461 (N4103, N4047, N4048);
nor NOR2_1462 (N4106, N1293_t0, N4049_t0);
nor NOR2_1463 (N4110, N4052_t0, N570_t0);
nor NOR2_1464 (N4114, N4055_t0, N618_t0);
nor NOR2_1465 (N4118, N4058_t0, N666_t0);
nor NOR2_1466 (N4122, N4061_t0, N714_t0);
nor NOR2_1467 (N4126, N4064_t0, N762_t0);
nor NOR2_1468 (N4130, N4067_t0, N810_t0);
nor NOR2_1469 (N4134, N4070_t0, N858_t0);
nor NOR2_1470 (N4138, N4019_t1, N4073_t0);
nor NOR2_1471 (N4139, N4073_t1, N906_t1);
nor NOR2_1472 (N4140, N3917_t2, N4073_t2);
nor NOR2_1473 (N4143, N4077, N4078);
nor NOR2_1474 (N4146, N4082_t0, N4079_t0);
nor NOR2_1475 (N4150, N4031_t1, N4085_t0);
nor NOR2_1476 (N4151, N4085_t1, N4028_t1);
nor NOR2_1477 (N4152, N4089, N4090);
nor NOR2_1478 (N4155, N4091_t0, N1101_t0);
nor NOR2_1479 (N4159, N4040_t1, N4094_t0);
nor NOR2_1480 (N4160, N4094_t1, N1149_t1);
nor NOR2_1481 (N4161, N3938_t2, N4094_t2);
nor NOR2_1482 (N4164, N4098, N4099);
nor NOR2_1483 (N4167, N4103_t0, N4100_t0);
nor NOR2_1484 (N4171, N1293_t1, N4106_t0);
nor NOR2_1485 (N4172, N4106_t1, N4049_t1);
nor NOR2_1486 (N4173, N4052_t1, N4110_t0);
nor NOR2_1487 (N4174, N4110_t1, N570_t1);
nor NOR2_1488 (N4175, N3947_t2, N4110_t2);
nor NOR2_1489 (N4178, N4055_t1, N4114_t0);
nor NOR2_1490 (N4179, N4114_t1, N618_t1);
nor NOR2_1491 (N4180, N3951_t2, N4114_t2);
nor NOR2_1492 (N4183, N4058_t1, N4118_t0);
nor NOR2_1493 (N4184, N4118_t1, N666_t1);
nor NOR2_1494 (N4185, N3955_t2, N4118_t2);
nor NOR2_1495 (N4188, N4061_t1, N4122_t0);
nor NOR2_1496 (N4189, N4122_t1, N714_t1);
nor NOR2_1497 (N4190, N3959_t2, N4122_t2);
nor NOR2_1498 (N4193, N4064_t1, N4126_t0);
nor NOR2_1499 (N4194, N4126_t1, N762_t1);
nor NOR2_1500 (N4195, N3963_t2, N4126_t2);
nor NOR2_1501 (N4198, N4067_t1, N4130_t0);
nor NOR2_1502 (N4199, N4130_t1, N810_t1);
nor NOR2_1503 (N4200, N3967_t2, N4130_t2);
nor NOR2_1504 (N4203, N4070_t1, N4134_t0);
nor NOR2_1505 (N4204, N4134_t1, N858_t1);
nor NOR2_1506 (N4205, N3971_t2, N4134_t2);
nor NOR2_1507 (N4208, N4138, N4139);
nor NOR2_1508 (N4211, N4143_t0, N4140_t0);
nor NOR2_1509 (N4215, N4082_t1, N4146_t0);
nor NOR2_1510 (N4216, N4146_t1, N4079_t1);
nor NOR2_1511 (N4217, N4150, N4151);
nor NOR2_1512 (N4220, N4152_t0, N1053_t0);
nor NOR2_1513 (N4224, N4091_t1, N4155_t0);
nor NOR2_1514 (N4225, N4155_t1, N1101_t1);
nor NOR2_1515 (N4226, N3992_t2, N4155_t2);
nor NOR2_1516 (N4229, N4159, N4160);
nor NOR2_1517 (N4232, N4164_t0, N4161_t0);
nor NOR2_1518 (N4236, N4103_t1, N4167_t0);
nor NOR2_1519 (N4237, N4167_t1, N4100_t1);
nor NOR2_1520 (N4238, N4171, N4172);
nor NOR2_1521 (N4241, N4173, N4174);
nor NOR2_1522 (N4242, N4178, N4179);
nor NOR2_1523 (N4245, N4183, N4184);
nor NOR2_1524 (N4248, N4188, N4189);
nor NOR2_1525 (N4251, N4193, N4194);
nor NOR2_1526 (N4254, N4198, N4199);
nor NOR2_1527 (N4257, N4203, N4204);
nor NOR2_1528 (N4260, N4208_t0, N4205_t0);
nor NOR2_1529 (N4264, N4143_t1, N4211_t0);
nor NOR2_1530 (N4265, N4211_t1, N4140_t1);
nor NOR2_1531 (N4266, N4215, N4216);
nor NOR2_1532 (N4269, N4217_t0, N1005_t0);
nor NOR2_1533 (N4273, N4152_t1, N4220_t0);
nor NOR2_1534 (N4274, N4220_t1, N1053_t1);
nor NOR2_1535 (N4275, N4034_t2, N4220_t2);
nor NOR2_1536 (N4278, N4224, N4225);
nor NOR2_1537 (N4281, N4229_t0, N4226_t0);
nor NOR2_1538 (N4285, N4164_t1, N4232_t0);
nor NOR2_1539 (N4286, N4232_t1, N4161_t1);
nor NOR2_1540 (N4287, N4236, N4237);
nor NOR2_1541 (N4290, N4238_t0, N1248_t0);
nor NOR2_1542 (N4294, N4242_t0, N4175_t0);
nor NOR2_1543 (N4298, N4245_t0, N4180_t0);
nor NOR2_1544 (N4302, N4248_t0, N4185_t0);
nor NOR2_1545 (N4306, N4251_t0, N4190_t0);
nor NOR2_1546 (N4310, N4254_t0, N4195_t0);
nor NOR2_1547 (N4314, N4257_t0, N4200_t0);
nor NOR2_1548 (N4318, N4208_t1, N4260_t0);
nor NOR2_1549 (N4319, N4260_t1, N4205_t1);
nor NOR2_1550 (N4320, N4264, N4265);
nor NOR2_1551 (N4323, N4266_t0, N957_t0);
nor NOR2_1552 (N4327, N4217_t1, N4269_t0);
nor NOR2_1553 (N4328, N4269_t1, N1005_t1);
nor NOR2_1554 (N4329, N4085_t2, N4269_t2);
nor NOR2_1555 (N4332, N4273, N4274);
nor NOR2_1556 (N4335, N4278_t0, N4275_t0);
nor NOR2_1557 (N4339, N4229_t1, N4281_t0);
nor NOR2_1558 (N4340, N4281_t1, N4226_t1);
nor NOR2_1559 (N4341, N4285, N4286);
nor NOR2_1560 (N4344, N4287_t0, N1200_t0);
nor NOR2_1561 (N4348, N4238_t1, N4290_t0);
nor NOR2_1562 (N4349, N4290_t1, N1248_t1);
nor NOR2_1563 (N4350, N4106_t2, N4290_t2);
nor NOR2_1564 (N4353, N4242_t1, N4294_t0);
nor NOR2_1565 (N4354, N4294_t1, N4175_t1);
nor NOR2_1566 (N4355, N4245_t1, N4298_t0);
nor NOR2_1567 (N4356, N4298_t1, N4180_t1);
nor NOR2_1568 (N4357, N4248_t1, N4302_t0);
nor NOR2_1569 (N4358, N4302_t1, N4185_t1);
nor NOR2_1570 (N4359, N4251_t1, N4306_t0);
nor NOR2_1571 (N4360, N4306_t1, N4190_t1);
nor NOR2_1572 (N4361, N4254_t1, N4310_t0);
nor NOR2_1573 (N4362, N4310_t1, N4195_t1);
nor NOR2_1574 (N4363, N4257_t1, N4314_t0);
nor NOR2_1575 (N4364, N4314_t1, N4200_t1);
nor NOR2_1576 (N4365, N4318, N4319);
nor NOR2_1577 (N4368, N4320_t0, N909_t0);
nor NOR2_1578 (N4372, N4266_t1, N4323_t0);
nor NOR2_1579 (N4373, N4323_t1, N957_t1);
nor NOR2_1580 (N4374, N4146_t2, N4323_t2);
nor NOR2_1581 (N4377, N4327, N4328);
nor NOR2_1582 (N4380, N4332_t0, N4329_t0);
nor NOR2_1583 (N4384, N4278_t1, N4335_t0);
nor NOR2_1584 (N4385, N4335_t1, N4275_t1);
nor NOR2_1585 (N4386, N4339, N4340);
nor NOR2_1586 (N4389, N4341_t0, N1152_t0);
nor NOR2_1587 (N4393, N4287_t1, N4344_t0);
nor NOR2_1588 (N4394, N4344_t1, N1200_t1);
nor NOR2_1589 (N4395, N4167_t2, N4344_t2);
nor NOR2_1590 (N4398, N4348, N4349);
nor NOR2_1591 (N4401, N1296_t0, N4350_t0);
nor NOR2_1592 (N4405, N4353, N4354);
nor NOR2_1593 (N4408, N4355, N4356);
nor NOR2_1594 (N4411, N4357, N4358);
nor NOR2_1595 (N4414, N4359, N4360);
nor NOR2_1596 (N4417, N4361, N4362);
nor NOR2_1597 (N4420, N4363, N4364);
nor NOR2_1598 (N4423, N4365_t0, N861_t0);
nor NOR2_1599 (N4427, N4320_t1, N4368_t0);
nor NOR2_1600 (N4428, N4368_t1, N909_t1);
nor NOR2_1601 (N4429, N4211_t2, N4368_t2);
nor NOR2_1602 (N4432, N4372, N4373);
nor NOR2_1603 (N4435, N4377_t0, N4374_t0);
nor NOR2_1604 (N4439, N4332_t1, N4380_t0);
nor NOR2_1605 (N4440, N4380_t1, N4329_t1);
nor NOR2_1606 (N4441, N4384, N4385);
nor NOR2_1607 (N4444, N4386_t0, N1104_t0);
nor NOR2_1608 (N4448, N4341_t1, N4389_t0);
nor NOR2_1609 (N4449, N4389_t1, N1152_t1);
nor NOR2_1610 (N4450, N4232_t2, N4389_t2);
nor NOR2_1611 (N4453, N4393, N4394);
nor NOR2_1612 (N4456, N4398_t0, N4395_t0);
nor NOR2_1613 (N4460, N1296_t1, N4401_t0);
nor NOR2_1614 (N4461, N4401_t1, N4350_t1);
nor NOR2_1615 (N4462, N4405_t0, N573_t0);
nor NOR2_1616 (N4466, N4408_t0, N621_t0);
nor NOR2_1617 (N4470, N4411_t0, N669_t0);
nor NOR2_1618 (N4474, N4414_t0, N717_t0);
nor NOR2_1619 (N4478, N4417_t0, N765_t0);
nor NOR2_1620 (N4482, N4420_t0, N813_t0);
nor NOR2_1621 (N4486, N4365_t1, N4423_t0);
nor NOR2_1622 (N4487, N4423_t1, N861_t1);
nor NOR2_1623 (N4488, N4260_t2, N4423_t2);
nor NOR2_1624 (N4491, N4427, N4428);
nor NOR2_1625 (N4494, N4432_t0, N4429_t0);
nor NOR2_1626 (N4498, N4377_t1, N4435_t0);
nor NOR2_1627 (N4499, N4435_t1, N4374_t1);
nor NOR2_1628 (N4500, N4439, N4440);
nor NOR2_1629 (N4503, N4441_t0, N1056_t0);
nor NOR2_1630 (N4507, N4386_t1, N4444_t0);
nor NOR2_1631 (N4508, N4444_t1, N1104_t1);
nor NOR2_1632 (N4509, N4281_t2, N4444_t2);
nor NOR2_1633 (N4512, N4448, N4449);
nor NOR2_1634 (N4515, N4453_t0, N4450_t0);
nor NOR2_1635 (N4519, N4398_t1, N4456_t0);
nor NOR2_1636 (N4520, N4456_t1, N4395_t1);
nor NOR2_1637 (N4521, N4460, N4461);
nor NOR2_1638 (N4524, N4405_t1, N4462_t0);
nor NOR2_1639 (N4525, N4462_t1, N573_t1);
nor NOR2_1640 (N4526, N4294_t2, N4462_t2);
nor NOR2_1641 (N4529, N4408_t1, N4466_t0);
nor NOR2_1642 (N4530, N4466_t1, N621_t1);
nor NOR2_1643 (N4531, N4298_t2, N4466_t2);
nor NOR2_1644 (N4534, N4411_t1, N4470_t0);
nor NOR2_1645 (N4535, N4470_t1, N669_t1);
nor NOR2_1646 (N4536, N4302_t2, N4470_t2);
nor NOR2_1647 (N4539, N4414_t1, N4474_t0);
nor NOR2_1648 (N4540, N4474_t1, N717_t1);
nor NOR2_1649 (N4541, N4306_t2, N4474_t2);
nor NOR2_1650 (N4544, N4417_t1, N4478_t0);
nor NOR2_1651 (N4545, N4478_t1, N765_t1);
nor NOR2_1652 (N4546, N4310_t2, N4478_t2);
nor NOR2_1653 (N4549, N4420_t1, N4482_t0);
nor NOR2_1654 (N4550, N4482_t1, N813_t1);
nor NOR2_1655 (N4551, N4314_t2, N4482_t2);
nor NOR2_1656 (N4554, N4486, N4487);
nor NOR2_1657 (N4557, N4491_t0, N4488_t0);
nor NOR2_1658 (N4561, N4432_t1, N4494_t0);
nor NOR2_1659 (N4562, N4494_t1, N4429_t1);
nor NOR2_1660 (N4563, N4498, N4499);
nor NOR2_1661 (N4566, N4500_t0, N1008_t0);
nor NOR2_1662 (N4570, N4441_t1, N4503_t0);
nor NOR2_1663 (N4571, N4503_t1, N1056_t1);
nor NOR2_1664 (N4572, N4335_t2, N4503_t2);
nor NOR2_1665 (N4575, N4507, N4508);
nor NOR2_1666 (N4578, N4512_t0, N4509_t0);
nor NOR2_1667 (N4582, N4453_t1, N4515_t0);
nor NOR2_1668 (N4583, N4515_t1, N4450_t1);
nor NOR2_1669 (N4584, N4519, N4520);
nor NOR2_1670 (N4587, N4521_t0, N1251_t0);
nor NOR2_1671 (N4591, N4524, N4525);
nor NOR2_1672 (N4592, N4529, N4530);
nor NOR2_1673 (N4595, N4534, N4535);
nor NOR2_1674 (N4598, N4539, N4540);
nor NOR2_1675 (N4601, N4544, N4545);
nor NOR2_1676 (N4604, N4549, N4550);
nor NOR2_1677 (N4607, N4554_t0, N4551_t0);
nor NOR2_1678 (N4611, N4491_t1, N4557_t0);
nor NOR2_1679 (N4612, N4557_t1, N4488_t1);
nor NOR2_1680 (N4613, N4561, N4562);
nor NOR2_1681 (N4616, N4563_t0, N960_t0);
nor NOR2_1682 (N4620, N4500_t1, N4566_t0);
nor NOR2_1683 (N4621, N4566_t1, N1008_t1);
nor NOR2_1684 (N4622, N4380_t2, N4566_t2);
nor NOR2_1685 (N4625, N4570, N4571);
nor NOR2_1686 (N4628, N4575_t0, N4572_t0);
nor NOR2_1687 (N4632, N4512_t1, N4578_t0);
nor NOR2_1688 (N4633, N4578_t1, N4509_t1);
nor NOR2_1689 (N4634, N4582, N4583);
nor NOR2_1690 (N4637, N4584_t0, N1203_t0);
nor NOR2_1691 (N4641, N4521_t1, N4587_t0);
nor NOR2_1692 (N4642, N4587_t1, N1251_t1);
nor NOR2_1693 (N4643, N4401_t2, N4587_t2);
nor NOR2_1694 (N4646, N4592_t0, N4526_t0);
nor NOR2_1695 (N4650, N4595_t0, N4531_t0);
nor NOR2_1696 (N4654, N4598_t0, N4536_t0);
nor NOR2_1697 (N4658, N4601_t0, N4541_t0);
nor NOR2_1698 (N4662, N4604_t0, N4546_t0);
nor NOR2_1699 (N4666, N4554_t1, N4607_t0);
nor NOR2_1700 (N4667, N4607_t1, N4551_t1);
nor NOR2_1701 (N4668, N4611, N4612);
nor NOR2_1702 (N4671, N4613_t0, N912_t0);
nor NOR2_1703 (N4675, N4563_t1, N4616_t0);
nor NOR2_1704 (N4676, N4616_t1, N960_t1);
nor NOR2_1705 (N4677, N4435_t2, N4616_t2);
nor NOR2_1706 (N4680, N4620, N4621);
nor NOR2_1707 (N4683, N4625_t0, N4622_t0);
nor NOR2_1708 (N4687, N4575_t1, N4628_t0);
nor NOR2_1709 (N4688, N4628_t1, N4572_t1);
nor NOR2_1710 (N4689, N4632, N4633);
nor NOR2_1711 (N4692, N4634_t0, N1155_t0);
nor NOR2_1712 (N4696, N4584_t1, N4637_t0);
nor NOR2_1713 (N4697, N4637_t1, N1203_t1);
nor NOR2_1714 (N4698, N4456_t2, N4637_t2);
nor NOR2_1715 (N4701, N4641, N4642);
nor NOR2_1716 (N4704, N1299_t0, N4643_t0);
nor NOR2_1717 (N4708, N4592_t1, N4646_t0);
nor NOR2_1718 (N4709, N4646_t1, N4526_t1);
nor NOR2_1719 (N4710, N4595_t1, N4650_t0);
nor NOR2_1720 (N4711, N4650_t1, N4531_t1);
nor NOR2_1721 (N4712, N4598_t1, N4654_t0);
nor NOR2_1722 (N4713, N4654_t1, N4536_t1);
nor NOR2_1723 (N4714, N4601_t1, N4658_t0);
nor NOR2_1724 (N4715, N4658_t1, N4541_t1);
nor NOR2_1725 (N4716, N4604_t1, N4662_t0);
nor NOR2_1726 (N4717, N4662_t1, N4546_t1);
nor NOR2_1727 (N4718, N4666, N4667);
nor NOR2_1728 (N4721, N4668_t0, N864_t0);
nor NOR2_1729 (N4725, N4613_t1, N4671_t0);
nor NOR2_1730 (N4726, N4671_t1, N912_t1);
nor NOR2_1731 (N4727, N4494_t2, N4671_t2);
nor NOR2_1732 (N4730, N4675, N4676);
nor NOR2_1733 (N4733, N4680_t0, N4677_t0);
nor NOR2_1734 (N4737, N4625_t1, N4683_t0);
nor NOR2_1735 (N4738, N4683_t1, N4622_t1);
nor NOR2_1736 (N4739, N4687, N4688);
nor NOR2_1737 (N4742, N4689_t0, N1107_t0);
nor NOR2_1738 (N4746, N4634_t1, N4692_t0);
nor NOR2_1739 (N4747, N4692_t1, N1155_t1);
nor NOR2_1740 (N4748, N4515_t2, N4692_t2);
nor NOR2_1741 (N4751, N4696, N4697);
nor NOR2_1742 (N4754, N4701_t0, N4698_t0);
nor NOR2_1743 (N4758, N1299_t1, N4704_t0);
nor NOR2_1744 (N4759, N4704_t1, N4643_t1);
nor NOR2_1745 (N4760, N4708, N4709);
nor NOR2_1746 (N4763, N4710, N4711);
nor NOR2_1747 (N4766, N4712, N4713);
nor NOR2_1748 (N4769, N4714, N4715);
nor NOR2_1749 (N4772, N4716, N4717);
nor NOR2_1750 (N4775, N4718_t0, N816_t0);
nor NOR2_1751 (N4779, N4668_t1, N4721_t0);
nor NOR2_1752 (N4780, N4721_t1, N864_t1);
nor NOR2_1753 (N4781, N4557_t2, N4721_t2);
nor NOR2_1754 (N4784, N4725, N4726);
nor NOR2_1755 (N4787, N4730_t0, N4727_t0);
nor NOR2_1756 (N4791, N4680_t1, N4733_t0);
nor NOR2_1757 (N4792, N4733_t1, N4677_t1);
nor NOR2_1758 (N4793, N4737, N4738);
nor NOR2_1759 (N4796, N4739_t0, N1059_t0);
nor NOR2_1760 (N4800, N4689_t1, N4742_t0);
nor NOR2_1761 (N4801, N4742_t1, N1107_t1);
nor NOR2_1762 (N4802, N4578_t2, N4742_t2);
nor NOR2_1763 (N4805, N4746, N4747);
nor NOR2_1764 (N4808, N4751_t0, N4748_t0);
nor NOR2_1765 (N4812, N4701_t1, N4754_t0);
nor NOR2_1766 (N4813, N4754_t1, N4698_t1);
nor NOR2_1767 (N4814, N4758, N4759);
nor NOR2_1768 (N4817, N4760_t0, N576_t0);
nor NOR2_1769 (N4821, N4763_t0, N624_t0);
nor NOR2_1770 (N4825, N4766_t0, N672_t0);
nor NOR2_1771 (N4829, N4769_t0, N720_t0);
nor NOR2_1772 (N4833, N4772_t0, N768_t0);
nor NOR2_1773 (N4837, N4718_t1, N4775_t0);
nor NOR2_1774 (N4838, N4775_t1, N816_t1);
nor NOR2_1775 (N4839, N4607_t2, N4775_t2);
nor NOR2_1776 (N4842, N4779, N4780);
nor NOR2_1777 (N4845, N4784_t0, N4781_t0);
nor NOR2_1778 (N4849, N4730_t1, N4787_t0);
nor NOR2_1779 (N4850, N4787_t1, N4727_t1);
nor NOR2_1780 (N4851, N4791, N4792);
nor NOR2_1781 (N4854, N4793_t0, N1011_t0);
nor NOR2_1782 (N4858, N4739_t1, N4796_t0);
nor NOR2_1783 (N4859, N4796_t1, N1059_t1);
nor NOR2_1784 (N4860, N4628_t2, N4796_t2);
nor NOR2_1785 (N4863, N4800, N4801);
nor NOR2_1786 (N4866, N4805_t0, N4802_t0);
nor NOR2_1787 (N4870, N4751_t1, N4808_t0);
nor NOR2_1788 (N4871, N4808_t1, N4748_t1);
nor NOR2_1789 (N4872, N4812, N4813);
nor NOR2_1790 (N4875, N4814_t0, N1254_t0);
nor NOR2_1791 (N4879, N4760_t1, N4817_t0);
nor NOR2_1792 (N4880, N4817_t1, N576_t1);
nor NOR2_1793 (N4881, N4646_t2, N4817_t2);
nor NOR2_1794 (N4884, N4763_t1, N4821_t0);
nor NOR2_1795 (N4885, N4821_t1, N624_t1);
nor NOR2_1796 (N4886, N4650_t2, N4821_t2);
nor NOR2_1797 (N4889, N4766_t1, N4825_t0);
nor NOR2_1798 (N4890, N4825_t1, N672_t1);
nor NOR2_1799 (N4891, N4654_t2, N4825_t2);
nor NOR2_1800 (N4894, N4769_t1, N4829_t0);
nor NOR2_1801 (N4895, N4829_t1, N720_t1);
nor NOR2_1802 (N4896, N4658_t2, N4829_t2);
nor NOR2_1803 (N4899, N4772_t1, N4833_t0);
nor NOR2_1804 (N4900, N4833_t1, N768_t1);
nor NOR2_1805 (N4901, N4662_t2, N4833_t2);
nor NOR2_1806 (N4904, N4837, N4838);
nor NOR2_1807 (N4907, N4842_t0, N4839_t0);
nor NOR2_1808 (N4911, N4784_t1, N4845_t0);
nor NOR2_1809 (N4912, N4845_t1, N4781_t1);
nor NOR2_1810 (N4913, N4849, N4850);
nor NOR2_1811 (N4916, N4851_t0, N963_t0);
nor NOR2_1812 (N4920, N4793_t1, N4854_t0);
nor NOR2_1813 (N4921, N4854_t1, N1011_t1);
nor NOR2_1814 (N4922, N4683_t2, N4854_t2);
nor NOR2_1815 (N4925, N4858, N4859);
nor NOR2_1816 (N4928, N4863_t0, N4860_t0);
nor NOR2_1817 (N4932, N4805_t1, N4866_t0);
nor NOR2_1818 (N4933, N4866_t1, N4802_t1);
nor NOR2_1819 (N4934, N4870, N4871);
nor NOR2_1820 (N4937, N4872_t0, N1206_t0);
nor NOR2_1821 (N4941, N4814_t1, N4875_t0);
nor NOR2_1822 (N4942, N4875_t1, N1254_t1);
nor NOR2_1823 (N4943, N4704_t2, N4875_t2);
nor NOR2_1824 (N4946, N4879, N4880);
nor NOR2_1825 (N4947, N4884, N4885);
nor NOR2_1826 (N4950, N4889, N4890);
nor NOR2_1827 (N4953, N4894, N4895);
nor NOR2_1828 (N4956, N4899, N4900);
nor NOR2_1829 (N4959, N4904_t0, N4901_t0);
nor NOR2_1830 (N4963, N4842_t1, N4907_t0);
nor NOR2_1831 (N4964, N4907_t1, N4839_t1);
nor NOR2_1832 (N4965, N4911, N4912);
nor NOR2_1833 (N4968, N4913_t0, N915_t0);
nor NOR2_1834 (N4972, N4851_t1, N4916_t0);
nor NOR2_1835 (N4973, N4916_t1, N963_t1);
nor NOR2_1836 (N4974, N4733_t2, N4916_t2);
nor NOR2_1837 (N4977, N4920, N4921);
nor NOR2_1838 (N4980, N4925_t0, N4922_t0);
nor NOR2_1839 (N4984, N4863_t1, N4928_t0);
nor NOR2_1840 (N4985, N4928_t1, N4860_t1);
nor NOR2_1841 (N4986, N4932, N4933);
nor NOR2_1842 (N4989, N4934_t0, N1158_t0);
nor NOR2_1843 (N4993, N4872_t1, N4937_t0);
nor NOR2_1844 (N4994, N4937_t1, N1206_t1);
nor NOR2_1845 (N4995, N4754_t2, N4937_t2);
nor NOR2_1846 (N4998, N4941, N4942);
nor NOR2_1847 (N5001, N1302_t0, N4943_t0);
nor NOR2_1848 (N5005, N4947_t0, N4881_t0);
nor NOR2_1849 (N5009, N4950_t0, N4886_t0);
nor NOR2_1850 (N5013, N4953_t0, N4891_t0);
nor NOR2_1851 (N5017, N4956_t0, N4896_t0);
nor NOR2_1852 (N5021, N4904_t1, N4959_t0);
nor NOR2_1853 (N5022, N4959_t1, N4901_t1);
nor NOR2_1854 (N5023, N4963, N4964);
nor NOR2_1855 (N5026, N4965_t0, N867_t0);
nor NOR2_1856 (N5030, N4913_t1, N4968_t0);
nor NOR2_1857 (N5031, N4968_t1, N915_t1);
nor NOR2_1858 (N5032, N4787_t2, N4968_t2);
nor NOR2_1859 (N5035, N4972, N4973);
nor NOR2_1860 (N5038, N4977_t0, N4974_t0);
nor NOR2_1861 (N5042, N4925_t1, N4980_t0);
nor NOR2_1862 (N5043, N4980_t1, N4922_t1);
nor NOR2_1863 (N5044, N4984, N4985);
nor NOR2_1864 (N5047, N4986_t0, N1110_t0);
nor NOR2_1865 (N5051, N4934_t1, N4989_t0);
nor NOR2_1866 (N5052, N4989_t1, N1158_t1);
nor NOR2_1867 (N5053, N4808_t2, N4989_t2);
nor NOR2_1868 (N5056, N4993, N4994);
nor NOR2_1869 (N5059, N4998_t0, N4995_t0);
nor NOR2_1870 (N5063, N1302_t1, N5001_t0);
nor NOR2_1871 (N5064, N5001_t1, N4943_t1);
nor NOR2_1872 (N5065, N4947_t1, N5005_t0);
nor NOR2_1873 (N5066, N5005_t1, N4881_t1);
nor NOR2_1874 (N5067, N4950_t1, N5009_t0);
nor NOR2_1875 (N5068, N5009_t1, N4886_t1);
nor NOR2_1876 (N5069, N4953_t1, N5013_t0);
nor NOR2_1877 (N5070, N5013_t1, N4891_t1);
nor NOR2_1878 (N5071, N4956_t1, N5017_t0);
nor NOR2_1879 (N5072, N5017_t1, N4896_t1);
nor NOR2_1880 (N5073, N5021, N5022);
nor NOR2_1881 (N5076, N5023_t0, N819_t0);
nor NOR2_1882 (N5080, N4965_t1, N5026_t0);
nor NOR2_1883 (N5081, N5026_t1, N867_t1);
nor NOR2_1884 (N5082, N4845_t2, N5026_t2);
nor NOR2_1885 (N5085, N5030, N5031);
nor NOR2_1886 (N5088, N5035_t0, N5032_t0);
nor NOR2_1887 (N5092, N4977_t1, N5038_t0);
nor NOR2_1888 (N5093, N5038_t1, N4974_t1);
nor NOR2_1889 (N5094, N5042, N5043);
nor NOR2_1890 (N5097, N5044_t0, N1062_t0);
nor NOR2_1891 (N5101, N4986_t1, N5047_t0);
nor NOR2_1892 (N5102, N5047_t1, N1110_t1);
nor NOR2_1893 (N5103, N4866_t2, N5047_t2);
nor NOR2_1894 (N5106, N5051, N5052);
nor NOR2_1895 (N5109, N5056_t0, N5053_t0);
nor NOR2_1896 (N5113, N4998_t1, N5059_t0);
nor NOR2_1897 (N5114, N5059_t1, N4995_t1);
nor NOR2_1898 (N5115, N5063, N5064);
nor NOR2_1899 (N5118, N5065, N5066);
nor NOR2_1900 (N5121, N5067, N5068);
nor NOR2_1901 (N5124, N5069, N5070);
nor NOR2_1902 (N5127, N5071, N5072);
nor NOR2_1903 (N5130, N5073_t0, N771_t0);
nor NOR2_1904 (N5134, N5023_t1, N5076_t0);
nor NOR2_1905 (N5135, N5076_t1, N819_t1);
nor NOR2_1906 (N5136, N4907_t2, N5076_t2);
nor NOR2_1907 (N5139, N5080, N5081);
nor NOR2_1908 (N5142, N5085_t0, N5082_t0);
nor NOR2_1909 (N5146, N5035_t1, N5088_t0);
nor NOR2_1910 (N5147, N5088_t1, N5032_t1);
nor NOR2_1911 (N5148, N5092, N5093);
nor NOR2_1912 (N5151, N5094_t0, N1014_t0);
nor NOR2_1913 (N5155, N5044_t1, N5097_t0);
nor NOR2_1914 (N5156, N5097_t1, N1062_t1);
nor NOR2_1915 (N5157, N4928_t2, N5097_t2);
nor NOR2_1916 (N5160, N5101, N5102);
nor NOR2_1917 (N5163, N5106_t0, N5103_t0);
nor NOR2_1918 (N5167, N5056_t1, N5109_t0);
nor NOR2_1919 (N5168, N5109_t1, N5053_t1);
nor NOR2_1920 (N5169, N5113, N5114);
nor NOR2_1921 (N5172, N5115_t0, N1257_t0);
nor NOR2_1922 (N5176, N5118_t0, N579_t0);
nor NOR2_1923 (N5180, N5121_t0, N627_t0);
nor NOR2_1924 (N5184, N5124_t0, N675_t0);
nor NOR2_1925 (N5188, N5127_t0, N723_t0);
nor NOR2_1926 (N5192, N5073_t1, N5130_t0);
nor NOR2_1927 (N5193, N5130_t1, N771_t1);
nor NOR2_1928 (N5194, N4959_t2, N5130_t2);
nor NOR2_1929 (N5197, N5134, N5135);
nor NOR2_1930 (N5200, N5139_t0, N5136_t0);
nor NOR2_1931 (N5204, N5085_t1, N5142_t0);
nor NOR2_1932 (N5205, N5142_t1, N5082_t1);
nor NOR2_1933 (N5206, N5146, N5147);
nor NOR2_1934 (N5209, N5148_t0, N966_t0);
nor NOR2_1935 (N5213, N5094_t1, N5151_t0);
nor NOR2_1936 (N5214, N5151_t1, N1014_t1);
nor NOR2_1937 (N5215, N4980_t2, N5151_t2);
nor NOR2_1938 (N5218, N5155, N5156);
nor NOR2_1939 (N5221, N5160_t0, N5157_t0);
nor NOR2_1940 (N5225, N5106_t1, N5163_t0);
nor NOR2_1941 (N5226, N5163_t1, N5103_t1);
nor NOR2_1942 (N5227, N5167, N5168);
nor NOR2_1943 (N5230, N5169_t0, N1209_t0);
nor NOR2_1944 (N5234, N5115_t1, N5172_t0);
nor NOR2_1945 (N5235, N5172_t1, N1257_t1);
nor NOR2_1946 (N5236, N5001_t2, N5172_t2);
nor NOR2_1947 (N5239, N5118_t1, N5176_t0);
nor NOR2_1948 (N5240, N5176_t1, N579_t1);
nor NOR2_1949 (N5241, N5005_t2, N5176_t2);
nor NOR2_1950 (N5244, N5121_t1, N5180_t0);
nor NOR2_1951 (N5245, N5180_t1, N627_t1);
nor NOR2_1952 (N5246, N5009_t2, N5180_t2);
nor NOR2_1953 (N5249, N5124_t1, N5184_t0);
nor NOR2_1954 (N5250, N5184_t1, N675_t1);
nor NOR2_1955 (N5251, N5013_t2, N5184_t2);
nor NOR2_1956 (N5254, N5127_t1, N5188_t0);
nor NOR2_1957 (N5255, N5188_t1, N723_t1);
nor NOR2_1958 (N5256, N5017_t2, N5188_t2);
nor NOR2_1959 (N5259, N5192, N5193);
nor NOR2_1960 (N5262, N5197_t0, N5194_t0);
nor NOR2_1961 (N5266, N5139_t1, N5200_t0);
nor NOR2_1962 (N5267, N5200_t1, N5136_t1);
nor NOR2_1963 (N5268, N5204, N5205);
nor NOR2_1964 (N5271, N5206_t0, N918_t0);
nor NOR2_1965 (N5275, N5148_t1, N5209_t0);
nor NOR2_1966 (N5276, N5209_t1, N966_t1);
nor NOR2_1967 (N5277, N5038_t2, N5209_t2);
nor NOR2_1968 (N5280, N5213, N5214);
nor NOR2_1969 (N5283, N5218_t0, N5215_t0);
nor NOR2_1970 (N5287, N5160_t1, N5221_t0);
nor NOR2_1971 (N5288, N5221_t1, N5157_t1);
nor NOR2_1972 (N5289, N5225, N5226);
nor NOR2_1973 (N5292, N5227_t0, N1161_t0);
nor NOR2_1974 (N5296, N5169_t1, N5230_t0);
nor NOR2_1975 (N5297, N5230_t1, N1209_t1);
nor NOR2_1976 (N5298, N5059_t2, N5230_t2);
nor NOR2_1977 (N5301, N5234, N5235);
nor NOR2_1978 (N5304, N1305_t0, N5236_t0);
nor NOR2_1979 (N5308, N5239, N5240);
nor NOR2_1980 (N5309, N5244, N5245);
nor NOR2_1981 (N5312, N5249, N5250);
nor NOR2_1982 (N5315, N5254, N5255);
nor NOR2_1983 (N5318, N5259_t0, N5256_t0);
nor NOR2_1984 (N5322, N5197_t1, N5262_t0);
nor NOR2_1985 (N5323, N5262_t1, N5194_t1);
nor NOR2_1986 (N5324, N5266, N5267);
nor NOR2_1987 (N5327, N5268_t0, N870_t0);
nor NOR2_1988 (N5331, N5206_t1, N5271_t0);
nor NOR2_1989 (N5332, N5271_t1, N918_t1);
nor NOR2_1990 (N5333, N5088_t2, N5271_t2);
nor NOR2_1991 (N5336, N5275, N5276);
nor NOR2_1992 (N5339, N5280_t0, N5277_t0);
nor NOR2_1993 (N5343, N5218_t1, N5283_t0);
nor NOR2_1994 (N5344, N5283_t1, N5215_t1);
nor NOR2_1995 (N5345, N5287, N5288);
nor NOR2_1996 (N5348, N5289_t0, N1113_t0);
nor NOR2_1997 (N5352, N5227_t1, N5292_t0);
nor NOR2_1998 (N5353, N5292_t1, N1161_t1);
nor NOR2_1999 (N5354, N5109_t2, N5292_t2);
nor NOR2_2000 (N5357, N5296, N5297);
nor NOR2_2001 (N5360, N5301_t0, N5298_t0);
nor NOR2_2002 (N5364, N1305_t1, N5304_t0);
nor NOR2_2003 (N5365, N5304_t1, N5236_t1);
nor NOR2_2004 (N5366, N5309_t0, N5241_t0);
nor NOR2_2005 (N5370, N5312_t0, N5246_t0);
nor NOR2_2006 (N5374, N5315_t0, N5251_t0);
nor NOR2_2007 (N5378, N5259_t1, N5318_t0);
nor NOR2_2008 (N5379, N5318_t1, N5256_t1);
nor NOR2_2009 (N5380, N5322, N5323);
nor NOR2_2010 (N5383, N5324_t0, N822_t0);
nor NOR2_2011 (N5387, N5268_t1, N5327_t0);
nor NOR2_2012 (N5388, N5327_t1, N870_t1);
nor NOR2_2013 (N5389, N5142_t2, N5327_t2);
nor NOR2_2014 (N5392, N5331, N5332);
nor NOR2_2015 (N5395, N5336_t0, N5333_t0);
nor NOR2_2016 (N5399, N5280_t1, N5339_t0);
nor NOR2_2017 (N5400, N5339_t1, N5277_t1);
nor NOR2_2018 (N5401, N5343, N5344);
nor NOR2_2019 (N5404, N5345_t0, N1065_t0);
nor NOR2_2020 (N5408, N5289_t1, N5348_t0);
nor NOR2_2021 (N5409, N5348_t1, N1113_t1);
nor NOR2_2022 (N5410, N5163_t2, N5348_t2);
nor NOR2_2023 (N5413, N5352, N5353);
nor NOR2_2024 (N5416, N5357_t0, N5354_t0);
nor NOR2_2025 (N5420, N5301_t1, N5360_t0);
nor NOR2_2026 (N5421, N5360_t1, N5298_t1);
nor NOR2_2027 (N5422, N5364, N5365);
nor NOR2_2028 (N5425, N5309_t1, N5366_t0);
nor NOR2_2029 (N5426, N5366_t1, N5241_t1);
nor NOR2_2030 (N5427, N5312_t1, N5370_t0);
nor NOR2_2031 (N5428, N5370_t1, N5246_t1);
nor NOR2_2032 (N5429, N5315_t1, N5374_t0);
nor NOR2_2033 (N5430, N5374_t1, N5251_t1);
nor NOR2_2034 (N5431, N5378, N5379);
nor NOR2_2035 (N5434, N5380_t0, N774_t0);
nor NOR2_2036 (N5438, N5324_t1, N5383_t0);
nor NOR2_2037 (N5439, N5383_t1, N822_t1);
nor NOR2_2038 (N5440, N5200_t2, N5383_t2);
nor NOR2_2039 (N5443, N5387, N5388);
nor NOR2_2040 (N5446, N5392_t0, N5389_t0);
nor NOR2_2041 (N5450, N5336_t1, N5395_t0);
nor NOR2_2042 (N5451, N5395_t1, N5333_t1);
nor NOR2_2043 (N5452, N5399, N5400);
nor NOR2_2044 (N5455, N5401_t0, N1017_t0);
nor NOR2_2045 (N5459, N5345_t1, N5404_t0);
nor NOR2_2046 (N5460, N5404_t1, N1065_t1);
nor NOR2_2047 (N5461, N5221_t2, N5404_t2);
nor NOR2_2048 (N5464, N5408, N5409);
nor NOR2_2049 (N5467, N5413_t0, N5410_t0);
nor NOR2_2050 (N5471, N5357_t1, N5416_t0);
nor NOR2_2051 (N5472, N5416_t1, N5354_t1);
nor NOR2_2052 (N5473, N5420, N5421);
nor NOR2_2053 (N5476, N5422_t0, N1260_t0);
nor NOR2_2054 (N5480, N5425, N5426);
nor NOR2_2055 (N5483, N5427, N5428);
nor NOR2_2056 (N5486, N5429, N5430);
nor NOR2_2057 (N5489, N5431_t0, N726_t0);
nor NOR2_2058 (N5493, N5380_t1, N5434_t0);
nor NOR2_2059 (N5494, N5434_t1, N774_t1);
nor NOR2_2060 (N5495, N5262_t2, N5434_t2);
nor NOR2_2061 (N5498, N5438, N5439);
nor NOR2_2062 (N5501, N5443_t0, N5440_t0);
nor NOR2_2063 (N5505, N5392_t1, N5446_t0);
nor NOR2_2064 (N5506, N5446_t1, N5389_t1);
nor NOR2_2065 (N5507, N5450, N5451);
nor NOR2_2066 (N5510, N5452_t0, N969_t0);
nor NOR2_2067 (N5514, N5401_t1, N5455_t0);
nor NOR2_2068 (N5515, N5455_t1, N1017_t1);
nor NOR2_2069 (N5516, N5283_t2, N5455_t2);
nor NOR2_2070 (N5519, N5459, N5460);
nor NOR2_2071 (N5522, N5464_t0, N5461_t0);
nor NOR2_2072 (N5526, N5413_t1, N5467_t0);
nor NOR2_2073 (N5527, N5467_t1, N5410_t1);
nor NOR2_2074 (N5528, N5471, N5472);
nor NOR2_2075 (N5531, N5473_t0, N1212_t0);
nor NOR2_2076 (N5535, N5422_t1, N5476_t0);
nor NOR2_2077 (N5536, N5476_t1, N1260_t1);
nor NOR2_2078 (N5537, N5304_t2, N5476_t2);
nor NOR2_2079 (N5540, N5480_t0, N582_t0);
nor NOR2_2080 (N5544, N5483_t0, N630_t0);
nor NOR2_2081 (N5548, N5486_t0, N678_t0);
nor NOR2_2082 (N5552, N5431_t1, N5489_t0);
nor NOR2_2083 (N5553, N5489_t1, N726_t1);
nor NOR2_2084 (N5554, N5318_t2, N5489_t2);
nor NOR2_2085 (N5557, N5493, N5494);
nor NOR2_2086 (N5560, N5498_t0, N5495_t0);
nor NOR2_2087 (N5564, N5443_t1, N5501_t0);
nor NOR2_2088 (N5565, N5501_t1, N5440_t1);
nor NOR2_2089 (N5566, N5505, N5506);
nor NOR2_2090 (N5569, N5507_t0, N921_t0);
nor NOR2_2091 (N5573, N5452_t1, N5510_t0);
nor NOR2_2092 (N5574, N5510_t1, N969_t1);
nor NOR2_2093 (N5575, N5339_t2, N5510_t2);
nor NOR2_2094 (N5578, N5514, N5515);
nor NOR2_2095 (N5581, N5519_t0, N5516_t0);
nor NOR2_2096 (N5585, N5464_t1, N5522_t0);
nor NOR2_2097 (N5586, N5522_t1, N5461_t1);
nor NOR2_2098 (N5587, N5526, N5527);
nor NOR2_2099 (N5590, N5528_t0, N1164_t0);
nor NOR2_2100 (N5594, N5473_t1, N5531_t0);
nor NOR2_2101 (N5595, N5531_t1, N1212_t1);
nor NOR2_2102 (N5596, N5360_t2, N5531_t2);
nor NOR2_2103 (N5599, N5535, N5536);
nor NOR2_2104 (N5602, N1308_t0, N5537_t0);
nor NOR2_2105 (N5606, N5480_t1, N5540_t0);
nor NOR2_2106 (N5607, N5540_t1, N582_t1);
nor NOR2_2107 (N5608, N5366_t2, N5540_t2);
nor NOR2_2108 (N5611, N5483_t1, N5544_t0);
nor NOR2_2109 (N5612, N5544_t1, N630_t1);
nor NOR2_2110 (N5613, N5370_t2, N5544_t2);
nor NOR2_2111 (N5616, N5486_t1, N5548_t0);
nor NOR2_2112 (N5617, N5548_t1, N678_t1);
nor NOR2_2113 (N5618, N5374_t2, N5548_t2);
nor NOR2_2114 (N5621, N5552, N5553);
nor NOR2_2115 (N5624, N5557_t0, N5554_t0);
nor NOR2_2116 (N5628, N5498_t1, N5560_t0);
nor NOR2_2117 (N5629, N5560_t1, N5495_t1);
nor NOR2_2118 (N5630, N5564, N5565);
nor NOR2_2119 (N5633, N5566_t0, N873_t0);
nor NOR2_2120 (N5637, N5507_t1, N5569_t0);
nor NOR2_2121 (N5638, N5569_t1, N921_t1);
nor NOR2_2122 (N5639, N5395_t2, N5569_t2);
nor NOR2_2123 (N5642, N5573, N5574);
nor NOR2_2124 (N5645, N5578_t0, N5575_t0);
nor NOR2_2125 (N5649, N5519_t1, N5581_t0);
nor NOR2_2126 (N5650, N5581_t1, N5516_t1);
nor NOR2_2127 (N5651, N5585, N5586);
nor NOR2_2128 (N5654, N5587_t0, N1116_t0);
nor NOR2_2129 (N5658, N5528_t1, N5590_t0);
nor NOR2_2130 (N5659, N5590_t1, N1164_t1);
nor NOR2_2131 (N5660, N5416_t2, N5590_t2);
nor NOR2_2132 (N5663, N5594, N5595);
nor NOR2_2133 (N5666, N5599_t0, N5596_t0);
nor NOR2_2134 (N5670, N1308_t1, N5602_t0);
nor NOR2_2135 (N5671, N5602_t1, N5537_t1);
nor NOR2_2136 (N5672, N5606, N5607);
nor NOR2_2137 (N5673, N5611, N5612);
nor NOR2_2138 (N5676, N5616, N5617);
nor NOR2_2139 (N5679, N5621_t0, N5618_t0);
nor NOR2_2140 (N5683, N5557_t1, N5624_t0);
nor NOR2_2141 (N5684, N5624_t1, N5554_t1);
nor NOR2_2142 (N5685, N5628, N5629);
nor NOR2_2143 (N5688, N5630_t0, N825_t0);
nor NOR2_2144 (N5692, N5566_t1, N5633_t0);
nor NOR2_2145 (N5693, N5633_t1, N873_t1);
nor NOR2_2146 (N5694, N5446_t2, N5633_t2);
nor NOR2_2147 (N5697, N5637, N5638);
nor NOR2_2148 (N5700, N5642_t0, N5639_t0);
nor NOR2_2149 (N5704, N5578_t1, N5645_t0);
nor NOR2_2150 (N5705, N5645_t1, N5575_t1);
nor NOR2_2151 (N5706, N5649, N5650);
nor NOR2_2152 (N5709, N5651_t0, N1068_t0);
nor NOR2_2153 (N5713, N5587_t1, N5654_t0);
nor NOR2_2154 (N5714, N5654_t1, N1116_t1);
nor NOR2_2155 (N5715, N5467_t2, N5654_t2);
nor NOR2_2156 (N5718, N5658, N5659);
nor NOR2_2157 (N5721, N5663_t0, N5660_t0);
nor NOR2_2158 (N5725, N5599_t1, N5666_t0);
nor NOR2_2159 (N5726, N5666_t1, N5596_t1);
nor NOR2_2160 (N5727, N5670, N5671);
nor NOR2_2161 (N5730, N5673_t0, N5608_t0);
nor NOR2_2162 (N5734, N5676_t0, N5613_t0);
nor NOR2_2163 (N5738, N5621_t1, N5679_t0);
nor NOR2_2164 (N5739, N5679_t1, N5618_t1);
nor NOR2_2165 (N5740, N5683, N5684);
nor NOR2_2166 (N5743, N5685_t0, N777_t0);
nor NOR2_2167 (N5747, N5630_t1, N5688_t0);
nor NOR2_2168 (N5748, N5688_t1, N825_t1);
nor NOR2_2169 (N5749, N5501_t2, N5688_t2);
nor NOR2_2170 (N5752, N5692, N5693);
nor NOR2_2171 (N5755, N5697_t0, N5694_t0);
nor NOR2_2172 (N5759, N5642_t1, N5700_t0);
nor NOR2_2173 (N5760, N5700_t1, N5639_t1);
nor NOR2_2174 (N5761, N5704, N5705);
nor NOR2_2175 (N5764, N5706_t0, N1020_t0);
nor NOR2_2176 (N5768, N5651_t1, N5709_t0);
nor NOR2_2177 (N5769, N5709_t1, N1068_t1);
nor NOR2_2178 (N5770, N5522_t2, N5709_t2);
nor NOR2_2179 (N5773, N5713, N5714);
nor NOR2_2180 (N5776, N5718_t0, N5715_t0);
nor NOR2_2181 (N5780, N5663_t1, N5721_t0);
nor NOR2_2182 (N5781, N5721_t1, N5660_t1);
nor NOR2_2183 (N5782, N5725, N5726);
nor NOR2_2184 (N5785, N5673_t1, N5730_t0);
nor NOR2_2185 (N5786, N5730_t1, N5608_t1);
nor NOR2_2186 (N5787, N5676_t1, N5734_t0);
nor NOR2_2187 (N5788, N5734_t1, N5613_t1);
nor NOR2_2188 (N5789, N5738, N5739);
nor NOR2_2189 (N5792, N5740_t0, N729_t0);
nor NOR2_2190 (N5796, N5685_t1, N5743_t0);
nor NOR2_2191 (N5797, N5743_t1, N777_t1);
nor NOR2_2192 (N5798, N5560_t2, N5743_t2);
nor NOR2_2193 (N5801, N5747, N5748);
nor NOR2_2194 (N5804, N5752_t0, N5749_t0);
nor NOR2_2195 (N5808, N5697_t1, N5755_t0);
nor NOR2_2196 (N5809, N5755_t1, N5694_t1);
nor NOR2_2197 (N5810, N5759, N5760);
nor NOR2_2198 (N5813, N5761_t0, N972_t0);
nor NOR2_2199 (N5817, N5706_t1, N5764_t0);
nor NOR2_2200 (N5818, N5764_t1, N1020_t1);
nor NOR2_2201 (N5819, N5581_t2, N5764_t2);
nor NOR2_2202 (N5822, N5768, N5769);
nor NOR2_2203 (N5825, N5773_t0, N5770_t0);
nor NOR2_2204 (N5829, N5718_t1, N5776_t0);
nor NOR2_2205 (N5830, N5776_t1, N5715_t1);
nor NOR2_2206 (N5831, N5780, N5781);
nor NOR2_2207 (N5834, N5785, N5786);
nor NOR2_2208 (N5837, N5787, N5788);
nor NOR2_2209 (N5840, N5789_t0, N681_t0);
nor NOR2_2210 (N5844, N5740_t1, N5792_t0);
nor NOR2_2211 (N5845, N5792_t1, N729_t1);
nor NOR2_2212 (N5846, N5624_t2, N5792_t2);
nor NOR2_2213 (N5849, N5796, N5797);
nor NOR2_2214 (N5852, N5801_t0, N5798_t0);
nor NOR2_2215 (N5856, N5752_t1, N5804_t0);
nor NOR2_2216 (N5857, N5804_t1, N5749_t1);
nor NOR2_2217 (N5858, N5808, N5809);
nor NOR2_2218 (N5861, N5810_t0, N924_t0);
nor NOR2_2219 (N5865, N5761_t1, N5813_t0);
nor NOR2_2220 (N5866, N5813_t1, N972_t1);
nor NOR2_2221 (N5867, N5645_t2, N5813_t2);
nor NOR2_2222 (N5870, N5817, N5818);
nor NOR2_2223 (N5873, N5822_t0, N5819_t0);
nor NOR2_2224 (N5877, N5773_t1, N5825_t0);
nor NOR2_2225 (N5878, N5825_t1, N5770_t1);
nor NOR2_2226 (N5879, N5829, N5830);
nor NOR2_2227 (N5882, N5834_t0, N585_t0);
nor NOR2_2228 (N5886, N5837_t0, N633_t0);
nor NOR2_2229 (N5890, N5789_t1, N5840_t0);
nor NOR2_2230 (N5891, N5840_t1, N681_t1);
nor NOR2_2231 (N5892, N5679_t2, N5840_t2);
nor NOR2_2232 (N5895, N5844, N5845);
nor NOR2_2233 (N5898, N5849_t0, N5846_t0);
nor NOR2_2234 (N5902, N5801_t1, N5852_t0);
nor NOR2_2235 (N5903, N5852_t1, N5798_t1);
nor NOR2_2236 (N5904, N5856, N5857);
nor NOR2_2237 (N5907, N5858_t0, N876_t0);
nor NOR2_2238 (N5911, N5810_t1, N5861_t0);
nor NOR2_2239 (N5912, N5861_t1, N924_t1);
nor NOR2_2240 (N5913, N5700_t2, N5861_t2);
nor NOR2_2241 (N5916, N5865, N5866);
nor NOR2_2242 (N5919, N5870_t0, N5867_t0);
nor NOR2_2243 (N5923, N5822_t1, N5873_t0);
nor NOR2_2244 (N5924, N5873_t1, N5819_t1);
nor NOR2_2245 (N5925, N5877, N5878);
nor NOR2_2246 (N5928, N5834_t1, N5882_t0);
nor NOR2_2247 (N5929, N5882_t1, N585_t1);
nor NOR2_2248 (N5930, N5730_t2, N5882_t2);
nor NOR2_2249 (N5933, N5837_t1, N5886_t0);
nor NOR2_2250 (N5934, N5886_t1, N633_t1);
nor NOR2_2251 (N5935, N5734_t2, N5886_t2);
nor NOR2_2252 (N5938, N5890, N5891);
nor NOR2_2253 (N5941, N5895_t0, N5892_t0);
nor NOR2_2254 (N5945, N5849_t1, N5898_t0);
nor NOR2_2255 (N5946, N5898_t1, N5846_t1);
nor NOR2_2256 (N5947, N5902, N5903);
nor NOR2_2257 (N5950, N5904_t0, N828_t0);
nor NOR2_2258 (N5954, N5858_t1, N5907_t0);
nor NOR2_2259 (N5955, N5907_t1, N876_t1);
nor NOR2_2260 (N5956, N5755_t2, N5907_t2);
nor NOR2_2261 (N5959, N5911, N5912);
nor NOR2_2262 (N5962, N5916_t0, N5913_t0);
nor NOR2_2263 (N5966, N5870_t1, N5919_t0);
nor NOR2_2264 (N5967, N5919_t1, N5867_t1);
nor NOR2_2265 (N5968, N5923, N5924);
nor NOR2_2266 (N5971, N5928, N5929);
nor NOR2_2267 (N5972, N5933, N5934);
nor NOR2_2268 (N5975, N5938_t0, N5935_t0);
nor NOR2_2269 (N5979, N5895_t1, N5941_t0);
nor NOR2_2270 (N5980, N5941_t1, N5892_t1);
nor NOR2_2271 (N5981, N5945, N5946);
nor NOR2_2272 (N5984, N5947_t0, N780_t0);
nor NOR2_2273 (N5988, N5904_t1, N5950_t0);
nor NOR2_2274 (N5989, N5950_t1, N828_t1);
nor NOR2_2275 (N5990, N5804_t2, N5950_t2);
nor NOR2_2276 (N5993, N5954, N5955);
nor NOR2_2277 (N5996, N5959_t0, N5956_t0);
nor NOR2_2278 (N6000, N5916_t1, N5962_t0);
nor NOR2_2279 (N6001, N5962_t1, N5913_t1);
nor NOR2_2280 (N6002, N5966, N5967);
nor NOR2_2281 (N6005, N5972_t0, N5930_t0);
nor NOR2_2282 (N6009, N5938_t1, N5975_t0);
nor NOR2_2283 (N6010, N5975_t1, N5935_t1);
nor NOR2_2284 (N6011, N5979, N5980);
nor NOR2_2285 (N6014, N5981_t0, N732_t0);
nor NOR2_2286 (N6018, N5947_t1, N5984_t0);
nor NOR2_2287 (N6019, N5984_t1, N780_t1);
nor NOR2_2288 (N6020, N5852_t2, N5984_t2);
nor NOR2_2289 (N6023, N5988, N5989);
nor NOR2_2290 (N6026, N5993_t0, N5990_t0);
nor NOR2_2291 (N6030, N5959_t1, N5996_t0);
nor NOR2_2292 (N6031, N5996_t1, N5956_t1);
nor NOR2_2293 (N6032, N6000, N6001);
nor NOR2_2294 (N6035, N5972_t1, N6005_t0);
nor NOR2_2295 (N6036, N6005_t1, N5930_t1);
nor NOR2_2296 (N6037, N6009, N6010);
nor NOR2_2297 (N6040, N6011_t0, N684_t0);
nor NOR2_2298 (N6044, N5981_t1, N6014_t0);
nor NOR2_2299 (N6045, N6014_t1, N732_t1);
nor NOR2_2300 (N6046, N5898_t2, N6014_t2);
nor NOR2_2301 (N6049, N6018, N6019);
nor NOR2_2302 (N6052, N6023_t0, N6020_t0);
nor NOR2_2303 (N6056, N5993_t1, N6026_t0);
nor NOR2_2304 (N6057, N6026_t1, N5990_t1);
nor NOR2_2305 (N6058, N6030, N6031);
nor NOR2_2306 (N6061, N6035, N6036);
nor NOR2_2307 (N6064, N6037_t0, N636_t0);
nor NOR2_2308 (N6068, N6011_t1, N6040_t0);
nor NOR2_2309 (N6069, N6040_t1, N684_t1);
nor NOR2_2310 (N6070, N5941_t2, N6040_t2);
nor NOR2_2311 (N6073, N6044, N6045);
nor NOR2_2312 (N6076, N6049_t0, N6046_t0);
nor NOR2_2313 (N6080, N6023_t1, N6052_t0);
nor NOR2_2314 (N6081, N6052_t1, N6020_t1);
nor NOR2_2315 (N6082, N6056, N6057);
nor NOR2_2316 (N6085, N6061_t0, N588_t0);
nor NOR2_2317 (N6089, N6037_t1, N6064_t0);
nor NOR2_2318 (N6090, N6064_t1, N636_t1);
nor NOR2_2319 (N6091, N5975_t2, N6064_t2);
nor NOR2_2320 (N6094, N6068, N6069);
nor NOR2_2321 (N6097, N6073_t0, N6070_t0);
nor NOR2_2322 (N6101, N6049_t1, N6076_t0);
nor NOR2_2323 (N6102, N6076_t1, N6046_t1);
nor NOR2_2324 (N6103, N6080, N6081);
nor NOR2_2325 (N6106, N6061_t1, N6085_t0);
nor NOR2_2326 (N6107, N6085_t1, N588_t1);
nor NOR2_2327 (N6108, N6005_t2, N6085_t2);
nor NOR2_2328 (N6111, N6089, N6090);
nor NOR2_2329 (N6114, N6094_t0, N6091_t0);
nor NOR2_2330 (N6118, N6073_t1, N6097_t0);
nor NOR2_2331 (N6119, N6097_t1, N6070_t1);
nor NOR2_2332 (N6120, N6101, N6102);
nor NOR2_2333 (N6123, N6106, N6107);
nor NOR2_2334 (N6124, N6111_t0, N6108_t0);
nor NOR2_2335 (N6128, N6094_t1, N6114_t0);
nor NOR2_2336 (N6129, N6114_t1, N6091_t1);
nor NOR2_2337 (N6130, N6118, N6119);
nor NOR2_2338 (N6133, N6111_t1, N6124_t0);
nor NOR2_2339 (N6134, N6124_t1, N6108_t1);
nor NOR2_2340 (N6135, N6128, N6129);
nor NOR2_2341 (N6138, N6133, N6134);
not NOT1_2342 (N6141, N6138_t0);
nor NOR2_2343 (N6145, N6138_t1, N6141_t0);
not NOT1_2344 (N6146, N6141_t1);
nor NOR2_2345 (N6147, N6124_t2, N6141_t2);
nor NOR2_2346 (N6150, N6145, N6146);
nor NOR2_2347 (N6151, N6135_t0, N6147_t0);
nor NOR2_2348 (N6155, N6135_t1, N6151_t0);
nor NOR2_2349 (N6156, N6151_t1, N6147_t1);
nor NOR2_2350 (N6157, N6114_t2, N6151_t2);
nor NOR2_2351 (N6160, N6155, N6156);
nor NOR2_2352 (N6161, N6130_t0, N6157_t0);
nor NOR2_2353 (N6165, N6130_t1, N6161_t0);
nor NOR2_2354 (N6166, N6161_t1, N6157_t1);
nor NOR2_2355 (N6167, N6097_t2, N6161_t2);
nor NOR2_2356 (N6170, N6165, N6166);
nor NOR2_2357 (N6171, N6120_t0, N6167_t0);
nor NOR2_2358 (N6175, N6120_t1, N6171_t0);
nor NOR2_2359 (N6176, N6171_t1, N6167_t1);
nor NOR2_2360 (N6177, N6076_t2, N6171_t2);
nor NOR2_2361 (N6180, N6175, N6176);
nor NOR2_2362 (N6181, N6103_t0, N6177_t0);
nor NOR2_2363 (N6185, N6103_t1, N6181_t0);
nor NOR2_2364 (N6186, N6181_t1, N6177_t1);
nor NOR2_2365 (N6187, N6052_t2, N6181_t2);
nor NOR2_2366 (N6190, N6185, N6186);
nor NOR2_2367 (N6191, N6082_t0, N6187_t0);
nor NOR2_2368 (N6195, N6082_t1, N6191_t0);
nor NOR2_2369 (N6196, N6191_t1, N6187_t1);
nor NOR2_2370 (N6197, N6026_t2, N6191_t2);
nor NOR2_2371 (N6200, N6195, N6196);
nor NOR2_2372 (N6201, N6058_t0, N6197_t0);
nor NOR2_2373 (N6205, N6058_t1, N6201_t0);
nor NOR2_2374 (N6206, N6201_t1, N6197_t1);
nor NOR2_2375 (N6207, N5996_t2, N6201_t2);
nor NOR2_2376 (N6210, N6205, N6206);
nor NOR2_2377 (N6211, N6032_t0, N6207_t0);
nor NOR2_2378 (N6215, N6032_t1, N6211_t0);
nor NOR2_2379 (N6216, N6211_t1, N6207_t1);
nor NOR2_2380 (N6217, N5962_t2, N6211_t2);
nor NOR2_2381 (N6220, N6215, N6216);
nor NOR2_2382 (N6221, N6002_t0, N6217_t0);
nor NOR2_2383 (N6225, N6002_t1, N6221_t0);
nor NOR2_2384 (N6226, N6221_t1, N6217_t1);
nor NOR2_2385 (N6227, N5919_t2, N6221_t2);
nor NOR2_2386 (N6230, N6225, N6226);
nor NOR2_2387 (N6231, N5968_t0, N6227_t0);
nor NOR2_2388 (N6235, N5968_t1, N6231_t0);
nor NOR2_2389 (N6236, N6231_t1, N6227_t1);
nor NOR2_2390 (N6237, N5873_t2, N6231_t2);
nor NOR2_2391 (N6240, N6235, N6236);
nor NOR2_2392 (N6241, N5925_t0, N6237_t0);
nor NOR2_2393 (N6245, N5925_t1, N6241_t0);
nor NOR2_2394 (N6246, N6241_t1, N6237_t1);
nor NOR2_2395 (N6247, N5825_t2, N6241_t2);
nor NOR2_2396 (N6250, N6245, N6246);
nor NOR2_2397 (N6251, N5879_t0, N6247_t0);
nor NOR2_2398 (N6255, N5879_t1, N6251_t0);
nor NOR2_2399 (N6256, N6251_t1, N6247_t1);
nor NOR2_2400 (N6257, N5776_t2, N6251_t2);
nor NOR2_2401 (N6260, N6255, N6256);
nor NOR2_2402 (N6261, N5831_t0, N6257_t0);
nor NOR2_2403 (N6265, N5831_t1, N6261_t0);
nor NOR2_2404 (N6266, N6261_t1, N6257_t1);
nor NOR2_2405 (N6267, N5721_t2, N6261_t2);
nor NOR2_2406 (N6270, N6265, N6266);
nor NOR2_2407 (N6271, N5782_t0, N6267_t0);
nor NOR2_2408 (N6275, N5782_t1, N6271_t0);
nor NOR2_2409 (N6276, N6271_t1, N6267_t1);
nor NOR2_2410 (N6277, N5666_t2, N6271_t2);
nor NOR2_2411 (N6280, N6275, N6276);
nor NOR2_2412 (N6281, N5727_t0, N6277_t0);
nor NOR2_2413 (N6285, N5727_t1, N6281_t0);
nor NOR2_2414 (N6286, N6281_t1, N6277_t1);
nor NOR2_2415 (N6287, N5602_t2, N6281_t2);
nor NOR2_2416 (N6288, N6285, N6286);

endmodule
