// Verilog
// c7552
// Ninputs 207
// Noutputs 108
// NtotalGates 3513
// BUFF1 535
// NOT1 876
// AND2 534
// AND4 64
// NAND2 1028
// NOR2 40
// OR2 180
// OR3 10
// AND5 32
// AND3 146
// OR5 24
// OR4 30
// NOR3 10
// NOR4 4

module c7552f (INC,END,clk,rst,N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
              N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
              N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
              N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
              N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
              N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
              N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
              N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
              N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
              N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
              N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
              N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
              N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
              N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
              N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
              N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
              N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
              N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
              N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
              N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
              N355,N358,N361,N364,N367,N382,N241_I,N387,N388,N478,
              N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,
              N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,
              N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,
              N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,
              N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,
              N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,
              N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,
              N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,N10716,N10717,
              N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,
              N10839,N10840,N10868,N10869,N10870,N10871,N10905,N10906,N10907,N10908,
              N11333,N11334,N11340,N11342,N241_O);

input N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
      N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
      N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
      N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
      N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
      N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
      N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
      N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
      N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
      N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
      N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
      N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
      N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
      N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
      N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
      N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
      N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
      N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
      N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
      N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
      N355,N358,N361,N364,N367,N382,N241_I;

output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,
       N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,
       N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,
       N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,
       N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,
       N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,
       N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,
       N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,
       N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,
       N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,
       N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;

wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,
     N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,
     N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,
     N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,
     N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,
     N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,
     N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,
     N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,
     N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,
     N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,
     N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,
     N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,
     N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,
     N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,
     N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,
     N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,
     N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,
     N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,
     N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,
     N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
     N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,
     N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,
     N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,
     N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
     N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,
     N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,
     N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
     N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
     N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
     N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,
     N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,
     N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,
     N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,
     N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,
     N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,
     N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
     N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,
     N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,
     N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,
     N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,
     N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,
     N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,
     N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
     N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
     N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,
     N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,
     N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,
     N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
     N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,
     N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,
     N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,
     N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,
     N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,
     N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,
     N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,
     N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,
     N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,
     N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
     N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,
     N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,
     N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,
     N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,
     N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,
     N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,
     N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,
     N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,
     N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,
     N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,
     N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,
     N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,
     N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,
     N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,
     N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,
     N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,
     N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,
     N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,
     N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,
     N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,
     N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,
     N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,
     N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,
     N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,
     N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,
     N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,
     N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,
     N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,
     N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,
     N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,
     N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
     N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
     N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,
     N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,
     N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
     N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
     N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,
     N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,
     N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,
     N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,
     N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,
     N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,
     N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
     N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,
     N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,
     N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,
     N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,
     N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,
     N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
     N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
     N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,
     N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,
     N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,
     N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,
     N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,
     N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,
     N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,
     N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,
     N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,
     N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,
     N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,
     N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,
     N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,
     N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,
     N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,
     N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
     N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,
     N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
     N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,
     N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,
     N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,
     N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,
     N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,
     N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,
     N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,
     N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,
     N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,
     N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,
     N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,
     N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,
     N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
     N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,
     N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,
     N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,
     N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,
     N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,
     N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,
     N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
     N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,
     N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,
     N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,
     N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,
     N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,
     N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,
     N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,
     N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,
     N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,
     N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,
     N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,
     N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,
     N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,
     N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,
     N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,
     N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,
     N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,
     N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,
     N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,
     N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
     N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,
     N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,
     N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,
     N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,
     N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,
     N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,
     N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,
     N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,
     N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,
     N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
     N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,
     N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,
     N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,
     N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,
     N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,
     N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
     N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,
     N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,
     N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,
     N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,
     N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,
     N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,
     N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,
     N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,
     N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,
     N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,
     N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,
     N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,
     N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,
     N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,
     N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,
     N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,
     N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,
     N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,
     N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,
     N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,
     N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,
     N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,
     N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,
     N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,
     N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,
     N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
     N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,
     N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,
     N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,
     N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,
     N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,
     N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,
     N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,
     N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,
     N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,
     N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,
     N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,
     N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,
     N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,
     N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,
     N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,
     N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,
     N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,
     N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,
     N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,
     N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,
     N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,
     N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,
     N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,
     N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,
     N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,
     N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,
     N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,
     N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,
     N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,
     N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,
     N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,
     N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
     N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,
     N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,
     N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,
     N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,
     N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,
     N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
     N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,
     N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,
     N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,
     N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,
     N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,
     N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,
     N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,
     N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,
     N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,
     N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,
     N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,
     N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,
     N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,
     N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,
     N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,
     N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,
     N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,
     N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
     N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,
     N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,
     N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,
     N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,
     N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,
     N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,
     N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,
     N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,
     N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,
     N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,
     N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,
     N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,
     N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,
     N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,
     N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,
     N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,
     N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,
     N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,
     N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,
     N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,
     N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,
     N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,
     N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,
     N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,
     N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,
     N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,
     N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,
     N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,
     N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,
     N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,
     N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,
     N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,
     N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,
     N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,
     N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,
     N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,
     N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
     N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,
     N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,
     N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,
     N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,
     N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,
     N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,
     N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,
     N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,
     N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,
     N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,
     N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,
     N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,
     N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,
     N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,
     N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,
     N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,
     N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,
     N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,
     N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,
     N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,
     N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,
     N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,
     N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,
     N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,
     N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,
     N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,
     N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
     N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,
     N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,
     N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,
     N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,
     N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,
     N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,
     N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,
     N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,
     N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,
     N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,
     N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,
     N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,
     N11336,N11337,N11338,N11339,N11341;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N53_t,N54_t,N55_t,N56_t,N57_t,N58_t,N59_t,N60_t,N61_t,N62_t,
     N63_t,N64_t,N65_t,N69_t,N73_t,N74_t,N75_t,N76_t,N77_t,N78_t,
     N79_t,N80_t,N81_t,N82_t,N83_t,N84_t,N85_t,N86_t,N87_t,N88_t,
     N109_t,N110_t,N111_t,N112_t,N113_t,N114_t,N133_t,N134_t,N150_t,N151_t,
     N152_t,N153_t,N154_t,N155_t,N156_t,N157_t,N158_t,N159_t,N160_t,N161_t,
     N162_t,N163_t,N164_t,N165_t,N166_t,N167_t,N168_t,N169_t,N170_t,N171_t,
     N172_t,N173_t,N174_t,N175_t,N176_t,N177_t,N178_t,N179_t,N180_t,N181_t,
     N182_t,N183_t,N184_t,N185_t,N186_t,N187_t,N188_t,N189_t,N190_t,N191_t,
     N192_t,N193_t,N194_t,N195_t,N196_t,N197_t,N198_t,N199_t,N200_t,N201_t,
     N202_t,N203_t,N204_t,N205_t,N206_t,N207_t,N208_t,N209_t,N210_t,N211_t,
     N212_t,N213_t,N214_t,N215_t,N216_t,N217_t,N218_t,N219_t,N220_t,N221_t,
     N222_t,N223_t,N224_t,N225_t,N226_t,N227_t,N228_t,N229_t,N230_t,N231_t,
     N232_t,N233_t,N234_t,N235_t,N236_t,N237_t,N238_t,N239_t,N240_t,N241_I_t;

     wire N1_t0,N1_t1,N1_t2,N248_t0,N248_t1,N254_t0,N254_t1,N257_t0,N257_t1,
     N260_t0,N260_t1,N263_t0,N263_t1,N263_t2,N267_t0,N267_t1,N267_t2,N274_t0,N274_t1,
     N280_t0,N280_t1,N283_t0,N283_t1,N286_t0,N286_t1,N289_t0,N289_t1,N289_t2,N293_t0,
     N293_t1,N296_t0,N296_t1,N299_t0,N299_t1,N299_t2,N303_t0,N303_t1,N303_t2,N307_t0,
     N307_t1,N310_t0,N310_t1,N313_t0,N313_t1,N316_t0,N316_t1,N319_t0,N319_t1,N322_t0,
     N322_t1,N325_t0,N325_t1,N328_t0,N328_t1,N331_t0,N331_t1,N334_t0,N334_t1,N337_t0,
     N337_t1,N343_t0,N343_t1,N346_t0,N346_t1,N349_t0,N349_t1,N352_t0,N352_t1,N355_t0,
     N355_t1,N358_t0,N358_t1,N361_t0,N361_t1,N364_t0,N364_t1,N15_t0,N15_t1,N5_t0,
     N5_t1,N5_t2,N38_t0,N38_t1,N12_t0,N12_t1,N9_t0,N9_t1,N245_t0,N245_t1,
     N251_t0,N251_t1,N106_t0,N106_t1,N18_t0,N18_t1,N18_t2,N18_t3,N382_t0,N382_t1,
     N382_t2,N382_t3,N271_t0,N271_t1,N277_t0,N277_t1,N367_t0,N367_t1,N367_t2,N367_t3,
     N367_t4,N367_t5,N367_t6,N367_t7,N367_t8,N367_t9,N367_t10,N367_t11,N367_t12,N367_t13,
     N340_t0,N340_t1,N528_t0,N528_t1,N578_t0,N578_t1,N575_t0,N575_t1,N494_t0,N494_t1,
     N590_t0,N590_t1,N657_t0,N657_t1,N469_t0,N469_t1,N596_t0,N596_t1,N242_t0,N242_t1,
     N593_t0,N593_t1,N625_t0,N625_t1,N871_t0,N871_t1,N628_t0,N628_t1,N628_t2,N682_t0,
     N682_t1,N682_t2,N682_t3,N682_t4,N632_t0,N632_t1,N632_t2,N676_t0,N676_t1,N676_t2,
     N676_t3,N676_t4,N700_t0,N700_t1,N700_t2,N700_t3,N614_t0,N614_t1,N614_t2,N614_t3,
     N614_t4,N614_t5,N614_t6,N614_t7,N614_t8,N614_t9,N689_t0,N689_t1,N689_t2,N689_t3,
     N689_t4,N695_t0,N695_t1,N695_t2,N695_t3,N750_t0,N750_t1,N750_t2,N750_t3,N666_t0,
     N666_t1,N666_t2,N666_t3,N666_t4,N660_t0,N660_t1,N660_t2,N660_t3,N660_t4,N651_t0,
     N651_t1,N651_t2,N651_t3,N651_t4,N644_t0,N644_t1,N644_t2,N644_t3,N644_t4,N644_t5,
     N609_t0,N609_t1,N609_t2,N609_t3,N604_t0,N604_t1,N604_t2,N604_t3,N742_t0,N742_t1,
     N742_t2,N742_t3,N742_t4,N599_t0,N599_t1,N599_t2,N599_t3,N727_t0,N727_t1,N727_t2,
     N727_t3,N727_t4,N721_t0,N721_t1,N721_t2,N721_t3,N721_t4,N715_t0,N715_t1,N715_t2,
     N715_t3,N715_t4,N734_t0,N734_t1,N734_t2,N734_t3,N734_t4,N734_t5,N734_t6,N708_t0,
     N708_t1,N708_t2,N708_t3,N708_t4,N708_t5,N806_t0,N806_t1,N806_t2,N806_t3,N806_t4,
     N800_t0,N800_t1,N800_t2,N800_t3,N800_t4,N794_t0,N794_t1,N794_t2,N794_t3,N794_t4,
     N786_t0,N786_t1,N786_t2,N786_t3,N786_t4,N786_t5,N786_t6,N780_t0,N780_t1,N780_t2,
     N780_t3,N780_t4,N774_t0,N774_t1,N774_t2,N774_t3,N774_t4,N768_t0,N768_t1,N768_t2,
     N768_t3,N768_t4,N762_t0,N762_t1,N762_t2,N762_t3,N762_t4,N636_t0,N636_t1,N636_t2,
     N636_t3,N865_t0,N865_t1,N865_t2,N865_t3,N865_t4,N859_t0,N859_t1,N859_t2,N859_t3,
     N859_t4,N853_t0,N853_t1,N853_t2,N853_t3,N853_t4,N845_t0,N845_t1,N845_t2,N845_t3,
     N845_t4,N845_t5,N845_t6,N839_t0,N839_t1,N839_t2,N839_t3,N839_t4,N833_t0,N833_t1,
     N833_t2,N833_t3,N833_t4,N827_t0,N827_t1,N827_t2,N827_t3,N827_t4,N821_t0,N821_t1,
     N821_t2,N821_t3,N821_t4,N814_t0,N814_t1,N814_t2,N814_t3,N814_t4,N814_t5,N1116_t0,
     N1116_t1,N957_t0,N957_t1,N957_t2,N957_t3,N957_t4,N957_t5,N1029_t0,N1029_t1,N1125_t0,
     N1125_t1,N1125_t2,N1125_t3,N1125_t4,N1125_t5,N1136_t0,N1136_t1,N1136_t2,N1136_t3,N1147_t0,
     N1147_t1,N1147_t2,N1147_t3,N1147_t4,N1147_t5,N1160_t0,N1160_t1,N1160_t2,N1160_t3,N1160_t4,
     N1160_t5,N1284_t0,N1284_t1,N1287_t0,N1287_t1,N1290_t0,N1290_t1,N1293_t0,N1293_t1,N1296_t0,
     N1296_t1,N1299_t0,N1299_t1,N1302_t0,N1302_t1,N1305_t0,N1305_t1,N1308_t0,N1308_t1,N1311_t0,
     N1311_t1,N1314_t0,N1314_t1,N1317_t0,N1317_t1,N1320_t0,N1320_t1,N1323_t0,N1323_t1,N1175_t0,
     N1175_t1,N1175_t2,N1175_t3,N1175_t4,N1175_t5,N1182_t0,N1182_t1,N1182_t2,N1182_t3,N1182_t4,
     N1182_t5,N1326_t0,N1326_t1,N1329_t0,N1329_t1,N1332_t0,N1332_t1,N1335_t0,N1335_t1,N1338_t0,
     N1338_t1,N1341_t0,N1341_t1,N1344_t0,N1344_t1,N1347_t0,N1347_t1,N1350_t0,N1350_t1,N1353_t0,
     N1353_t1,N1356_t0,N1356_t1,N1359_t0,N1359_t1,N1362_t0,N1362_t1,N1365_t0,N1365_t1,N1368_t0,
     N1368_t1,N1371_t0,N1371_t1,N1374_t0,N1374_t1,N1377_t0,N1377_t1,N1199_t0,N1199_t1,N1194_t0,
     N1194_t1,N1194_t2,N1194_t3,N1211_t0,N1211_t1,N1211_t2,N1211_t3,N1211_t4,N1211_t5,N44_t0,
     N44_t1,N41_t0,N41_t1,N29_t0,N29_t1,N26_t0,N26_t1,N23_t0,N23_t1,N1380_t0,
     N1380_t1,N1383_t0,N1383_t1,N1386_t0,N1386_t1,N1389_t0,N1389_t1,N1392_t0,N1392_t1,N1395_t0,
     N1395_t1,N1398_t0,N1398_t1,N1401_t0,N1401_t1,N1404_t0,N1404_t1,N1407_t0,N1407_t1,N1410_t0,
     N1410_t1,N1413_t0,N1413_t1,N1416_t0,N1416_t1,N1419_t0,N1419_t1,N1422_t0,N1422_t1,N1425_t0,
     N1425_t1,N1233_t0,N1233_t1,N1233_t2,N1233_t3,N1233_t4,N1233_t5,N1244_t0,N1244_t1,N1244_t2,
     N1244_t3,N1428_t0,N1428_t1,N1222_t0,N1222_t1,N1431_t0,N1431_t1,N1434_t0,N1434_t1,N1437_t0,
     N1437_t1,N1440_t0,N1440_t1,N1443_t0,N1443_t1,N1446_t0,N1446_t1,N1449_t0,N1449_t1,N1452_t0,
     N1452_t1,N1455_t0,N1455_t1,N1458_t0,N1458_t1,N1249_t0,N1249_t1,N1249_t2,N1249_t3,N1249_t4,
     N1249_t5,N1256_t0,N1256_t1,N1256_t2,N1256_t3,N1256_t4,N1256_t5,N1263_t0,N1263_t1,N1263_t2,
     N1263_t3,N1263_t4,N1263_t5,N47_t0,N47_t1,N35_t0,N35_t1,N32_t0,N32_t1,N50_t0,
     N50_t1,N66_t0,N66_t1,N1461_t0,N1461_t1,N1464_t0,N1464_t1,N1467_t0,N1467_t1,N1470_t0,
     N1470_t1,N1473_t0,N1473_t1,N1476_t0,N1476_t1,N1479_t0,N1479_t1,N1482_t0,N1482_t1,N1485_t0,
     N1485_t1,N1206_t0,N1206_t1,N1206_t2,N1206_t3,N1270_t0,N1270_t1,N1270_t2,N1270_t3,N1270_t4,
     N1270_t5,N1277_t0,N1277_t1,N1277_t2,N1277_t3,N1277_t4,N1277_t5,N1189_t0,N1189_t1,N1189_t2,
     N1189_t3,N1703_t0,N1703_t1,N1713_t0,N1713_t1,N1721_t0,N1721_t1,N1758_t0,N1758_t1,N1708_t0,
     N1708_t1,N1537_t0,N1537_t1,N1537_t2,N1537_t3,N1537_t4,N1551_t0,N1551_t1,N1783_t0,N1783_t1,
     N1783_t2,N1783_t3,N1783_t4,N1789_t0,N1789_t1,N1789_t2,N1799_t0,N1799_t1,N1799_t2,N1799_t3,
     N1799_t4,N1805_t0,N1805_t1,N1805_t2,N1805_t3,N1805_t4,N2074_t0,N2074_t1,N2081_t0,N2081_t1,
     N141_t0,N141_t1,N1845_t0,N1845_t1,N1845_t2,N1845_t3,N1845_t4,N147_t0,N147_t1,N138_t0,
     N138_t1,N144_t0,N144_t1,N135_t0,N135_t1,N1851_t0,N1851_t1,N1851_t2,N1851_t3,N1851_t4,
     N1885_t0,N1885_t1,N1885_t2,N1885_t3,N1885_t4,N1885_t5,N1892_t0,N1892_t1,N1892_t2,N1892_t3,
     N1892_t4,N1892_t5,N103_t0,N103_t1,N130_t0,N130_t1,N127_t0,N127_t1,N124_t0,N124_t1,
     N100_t0,N100_t1,N1899_t0,N1899_t1,N1899_t2,N1899_t3,N1899_t4,N1899_t5,N1906_t0,N1906_t1,
     N1906_t2,N1906_t3,N1906_t4,N1906_t5,N115_t0,N115_t1,N118_t0,N118_t1,N97_t0,N97_t1,
     N94_t0,N94_t1,N121_t0,N121_t1,N1919_t0,N1919_t1,N1919_t2,N1919_t3,N1919_t4,N1919_t5,
     N1913_t0,N1913_t1,N1913_t2,N1913_t3,N1913_t4,N1947_t0,N1947_t1,N1947_t2,N1947_t3,N1947_t4,
     N1953_t0,N1953_t1,N1953_t2,N2086_t0,N2086_t1,N1977_t0,N1977_t1,N1977_t2,N1977_t3,N1977_t4,
     N1983_t0,N1983_t1,N1983_t2,N1983_t3,N1983_t4,N759_t0,N759_t1,N70_t0,N70_t1,N2003_t0,
     N2003_t1,N2003_t2,N2003_t3,N2003_t4,N2003_t5,N1997_t0,N1997_t1,N1997_t2,N1997_t3,N1997_t4,
     N2024_t0,N2024_t1,N2024_t2,N2024_t3,N2024_t4,N2024_t5,N2031_t0,N2031_t1,N2031_t2,N2031_t3,
     N2031_t4,N2031_t5,N2038_t0,N2038_t1,N2038_t2,N2038_t3,N2038_t4,N2038_t5,N2045_t0,N2045_t1,
     N2045_t2,N2045_t3,N2045_t4,N2045_t5,N2052_t0,N2052_t1,N2052_t2,N2052_t3,N2052_t4,N2058_t0,
     N2058_t1,N2058_t2,N2058_t3,N2058_t4,N1119_t0,N1119_t1,N1119_t2,N1119_t3,N1119_t4,N1132_t0,
     N1132_t1,N1132_t2,N1141_t0,N1141_t1,N1141_t2,N1141_t3,N1141_t4,N1154_t0,N1154_t1,N1154_t2,
     N1154_t3,N1154_t4,N2235_t0,N2235_t1,N1227_t0,N1227_t1,N1227_t2,N1227_t3,N1227_t4,N1240_t0,
     N1240_t1,N1240_t2,N2231_t0,N2231_t1,N2257_t0,N2257_t1,N2257_t2,N2257_t3,N2257_t4,N2257_t5,
     N2257_t6,N2257_t7,N2257_t8,N2269_t0,N2269_t1,N2269_t2,N2269_t3,N2287_t0,N2287_t1,N2287_t2,
     N2287_t3,N2287_t4,N2293_t0,N2293_t1,N2293_t2,N2293_t3,N2293_t4,N2309_t0,N2309_t1,N2309_t2,
     N2309_t3,N2309_t4,N2315_t0,N2315_t1,N2315_t2,N2315_t3,N2315_t4,N2331_t0,N2331_t1,N2331_t2,
     N2331_t3,N2331_t4,N2368_t0,N2368_t1,N2368_t2,N2368_t3,N2368_t4,N2384_t0,N2384_t1,N2384_t2,
     N2384_t3,N2384_t4,N2390_t0,N2390_t1,N2390_t2,N2390_t3,N2390_t4,N2406_t0,N2406_t1,N2406_t2,
     N2406_t3,N2406_t4,N2412_t0,N2412_t1,N2412_t2,N2412_t3,N2412_t4,N2644_t0,N2644_t1,N2644_t2,
     N2644_t3,N2644_t4,N2638_t0,N2638_t1,N2638_t2,N2638_t3,N2638_t4,N2632_t0,N2632_t1,N2632_t2,
     N2632_t3,N2632_t4,N2626_t0,N2626_t1,N2626_t2,N2626_t3,N2626_t4,N2619_t0,N2619_t1,N2619_t2,
     N2619_t3,N2619_t4,N2619_t5,N2523_t0,N2523_t1,N2523_t2,N2523_t3,N2523_t4,N1167_t0,N1167_t1,
     N1167_t2,N1167_t3,N2533_t0,N2533_t1,N2533_t2,N2778_t0,N2778_t1,N2508_t0,N2508_t1,N2508_t2,
     N2508_t3,N2508_t4,N2502_t0,N2502_t1,N2502_t2,N2502_t3,N2502_t4,N2496_t0,N2496_t1,N2496_t2,
     N2496_t3,N2496_t4,N2488_t0,N2488_t1,N2488_t2,N2488_t3,N2488_t4,N2488_t5,N2488_t6,N2482_t0,
     N2482_t1,N2482_t2,N2482_t3,N2482_t4,N2573_t0,N2573_t1,N2573_t2,N2573_t3,N2573_t4,N2567_t0,
     N2567_t1,N2567_t2,N2567_t3,N2567_t4,N2561_t0,N2561_t1,N2561_t2,N2561_t3,N2561_t4,N2554_t0,
     N2554_t1,N2554_t2,N2554_t3,N2554_t4,N2554_t5,N2761_t0,N2761_t1,N2761_t2,N2478_t0,N2478_t1,
     N2478_t2,N2757_t0,N2757_t1,N2757_t2,N2474_t0,N2474_t1,N2474_t2,N2753_t0,N2753_t1,N2753_t2,
     N2470_t0,N2470_t1,N2470_t2,N2749_t0,N2749_t1,N2749_t2,N2466_t0,N2466_t1,N2466_t2,N2745_t0,
     N2745_t1,N2745_t2,N2462_t0,N2462_t1,N2462_t2,N2741_t0,N2741_t1,N2741_t2,N2550_t0,N2550_t1,
     N2550_t2,N2737_t0,N2737_t1,N2737_t2,N2546_t0,N2546_t1,N2546_t2,N2733_t0,N2733_t1,N2733_t2,
     N2542_t0,N2542_t1,N2542_t2,N2729_t0,N2729_t1,N2729_t2,N2538_t0,N2538_t1,N2538_t2,N2670_t0,
     N2670_t1,N2670_t2,N2458_t0,N2458_t1,N2458_t2,N2666_t0,N2666_t1,N2666_t2,N2454_t0,N2454_t1,
     N2454_t2,N2662_t0,N2662_t1,N2662_t2,N2450_t0,N2450_t1,N2450_t2,N2658_t0,N2658_t1,N2658_t2,
     N2446_t0,N2446_t1,N2446_t2,N2654_t0,N2654_t1,N2654_t2,N2442_t0,N2442_t1,N2442_t2,N2650_t0,
     N2650_t1,N2781_t0,N2781_t1,N2604_t0,N2604_t1,N2790_t0,N2790_t1,N2793_t0,N2793_t1,N2796_t0,
     N2796_t1,N2766_t0,N2766_t1,N2769_t0,N2769_t1,N2772_t0,N2772_t1,N2775_t0,N2775_t1,N2674_t0,
     N2674_t1,N2674_t2,N2674_t3,N2674_t4,N2704_t0,N2704_t1,N2704_t2,N2700_t0,N2700_t1,N2700_t2,
     N2696_t0,N2696_t1,N2696_t2,N2688_t0,N2688_t1,N2688_t2,N2692_t0,N2692_t1,N2692_t2,N2784_t0,
     N2784_t1,N2787_t0,N2787_t1,N2611_t0,N2611_t1,N2611_t2,N2607_t0,N2607_t1,N2607_t2,N2615_t0,
     N2615_t1,N2615_t2,N2680_t0,N2680_t1,N3067_t0,N3067_t1,N3070_t0,N3070_t1,N3073_t0,N3073_t1,
     N3080_t0,N3080_t1,N3061_t0,N3061_t1,N3064_t0,N3064_t1,N3487_t0,N3487_t1,N3490_t0,N3490_t1,
     N3493_t0,N3493_t1,N3496_t0,N3496_t1,N3499_t0,N3499_t1,N3122_t0,N3122_t1,N3122_t2,N3126_t0,
     N3126_t1,N3126_t2,N3518_t0,N3518_t1,N3521_t0,N3521_t1,N3524_t0,N3524_t1,N3527_t0,N3527_t1,
     N3530_t0,N3530_t1,N3155_t0,N3155_t1,N3155_t2,N3159_t0,N3159_t1,N3159_t2,N3535_t0,N3535_t1,
     N3539_t0,N3539_t1,N3542_t0,N3542_t1,N3545_t0,N3545_t1,N3548_t0,N3548_t1,N3553_t0,N3553_t1,
     N3557_t0,N3557_t1,N3560_t0,N3560_t1,N3563_t0,N3563_t1,N3566_t0,N3566_t1,N3571_t0,N3571_t1,
     N3574_t0,N3574_t1,N3577_t0,N3577_t1,N3580_t0,N3580_t1,N3583_t0,N3583_t1,N3598_t0,N3598_t1,
     N3601_t0,N3601_t1,N3604_t0,N3604_t1,N3607_t0,N3607_t1,N3610_t0,N3610_t1,N3613_t0,N3613_t1,
     N3616_t0,N3616_t1,N3619_t0,N3619_t1,N3622_t0,N3622_t1,N3631_t0,N3631_t1,N3634_t0,N3634_t1,
     N3637_t0,N3637_t1,N3640_t0,N3640_t1,N3643_t0,N3643_t1,N3646_t0,N3646_t1,N3649_t0,N3649_t1,
     N3652_t0,N3652_t1,N3655_t0,N3655_t1,N3658_t0,N3658_t1,N3293_t0,N3293_t1,N3293_t2,N3293_t3,
     N3293_t4,N3287_t0,N3287_t1,N3287_t2,N3287_t3,N3287_t4,N3281_t0,N3281_t1,N3281_t2,N3281_t3,
     N3281_t4,N3273_t0,N3273_t1,N3273_t2,N3273_t3,N3273_t4,N3273_t5,N3273_t6,N3267_t0,N3267_t1,
     N3267_t2,N3267_t3,N3267_t4,N3355_t0,N3355_t1,N3355_t2,N3355_t3,N3355_t4,N3349_t0,N3349_t1,
     N3349_t2,N3349_t3,N3349_t4,N3343_t0,N3343_t1,N3343_t2,N3343_t3,N3343_t4,N3661_t0,N3661_t1,
     N3664_t0,N3664_t1,N3667_t0,N3667_t1,N3670_t0,N3670_t1,N3673_t0,N3673_t1,N3676_t0,N3676_t1,
     N3679_t0,N3679_t1,N3682_t0,N3682_t1,N3685_t0,N3685_t1,N3688_t0,N3688_t1,N3691_t0,N3691_t1,
     N3694_t0,N3694_t1,N3697_t0,N3697_t1,N3700_t0,N3700_t1,N3703_t0,N3703_t1,N3706_t0,N3706_t1,
     N3709_t0,N3709_t1,N3712_t0,N3712_t1,N3715_t0,N3715_t1,N3718_t0,N3718_t1,N3721_t0,N3721_t1,
     N3448_t0,N3448_t1,N3448_t2,N3724_t0,N3724_t1,N3444_t0,N3444_t1,N3444_t2,N3727_t0,N3727_t1,
     N3440_t0,N3440_t1,N3440_t2,N3436_t0,N3436_t1,N3436_t2,N3730_t0,N3730_t1,N3432_t0,N3432_t1,
     N3432_t2,N3428_t0,N3428_t1,N3428_t2,N3311_t0,N3311_t1,N3311_t2,N3424_t0,N3424_t1,N3424_t2,
     N3307_t0,N3307_t1,N3307_t2,N3420_t0,N3420_t1,N3420_t2,N3303_t0,N3303_t1,N3303_t2,N3416_t0,
     N3416_t1,N3416_t2,N3299_t0,N3299_t1,N3299_t2,N3733_t0,N3733_t1,N3736_t0,N3736_t1,N3739_t0,
     N3739_t1,N3742_t0,N3742_t1,N3745_t0,N3745_t1,N3748_t0,N3748_t1,N3751_t0,N3751_t1,N3754_t0,
     N3754_t1,N3757_t0,N3757_t1,N3760_t0,N3760_t1,N3763_t0,N3763_t1,N3375_t0,N3375_t1,N3375_t2,
     N3410_t0,N3410_t1,N3410_t2,N3410_t3,N3410_t4,N3404_t0,N3404_t1,N3404_t2,N3404_t3,N3404_t4,
     N3398_t0,N3398_t1,N3398_t2,N3398_t3,N3398_t4,N3390_t0,N3390_t1,N3390_t2,N3390_t3,N3390_t4,
     N3390_t5,N3390_t6,N3384_t0,N3384_t1,N3384_t2,N3384_t3,N3384_t4,N3334_t0,N3334_t1,N3334_t2,
     N3334_t3,N3334_t4,N3328_t0,N3328_t1,N3328_t2,N3328_t3,N3328_t4,N3322_t0,N3322_t1,N3322_t2,
     N3322_t3,N3322_t4,N3315_t0,N3315_t1,N3315_t2,N3315_t3,N3315_t4,N3315_t5,N3766_t0,N3766_t1,
     N3769_t0,N3769_t1,N3772_t0,N3772_t1,N3775_t0,N3775_t1,N3778_t0,N3778_t1,N3783_t0,N3783_t1,
     N3786_t0,N3786_t1,N3789_t0,N3789_t1,N3792_t0,N3792_t1,N3807_t0,N3807_t1,N3810_t0,N3810_t1,
     N3813_t0,N3813_t1,N3816_t0,N3816_t1,N3819_t0,N3819_t1,N3822_t0,N3822_t1,N3825_t0,N3825_t1,
     N3828_t0,N3828_t1,N3831_t0,N3831_t1,N3482_t0,N3482_t1,N3482_t2,N3263_t0,N3263_t1,N3263_t2,
     N3478_t0,N3478_t1,N3478_t2,N3259_t0,N3259_t1,N3259_t2,N3474_t0,N3474_t1,N3474_t2,N3255_t0,
     N3255_t1,N3255_t2,N3470_t0,N3470_t1,N3470_t2,N3251_t0,N3251_t1,N3251_t2,N3466_t0,N3466_t1,
     N3466_t2,N3247_t0,N3247_t1,N3247_t2,N3846_t0,N3846_t1,N3462_t0,N3462_t1,N3462_t2,N3849_t0,
     N3849_t1,N3458_t0,N3458_t1,N3458_t2,N3852_t0,N3852_t1,N3454_t0,N3454_t1,N3454_t2,N3381_t0,
     N3381_t1,N3855_t0,N3855_t1,N3340_t0,N3340_t1,N3858_t0,N3858_t1,N3861_t0,N3861_t1,N3864_t0,
     N3864_t1,N3867_t0,N3867_t1,N3870_t0,N3870_t1,N3885_t0,N3885_t1,N3888_t0,N3888_t1,N3891_t0,
     N3891_t1,N3131_t0,N3131_t1,N3502_t0,N3502_t1,N3507_t0,N3507_t1,N3510_t0,N3510_t1,N3515_t0,
     N3515_t1,N3114_t0,N3114_t1,N3114_t2,N3114_t3,N3114_t4,N3114_t5,N3114_t6,N3586_t0,N3586_t1,
     N3589_t0,N3589_t1,N3592_t0,N3592_t1,N3595_t0,N3595_t1,N3625_t0,N3625_t1,N3178_t0,N3178_t1,
     N3178_t2,N3178_t3,N3178_t4,N3628_t0,N3628_t1,N3202_t0,N3202_t1,N3202_t2,N3202_t3,N3202_t4,
     N3202_t5,N3202_t6,N3221_t0,N3221_t1,N3221_t2,N3221_t3,N3221_t4,N3221_t5,N3795_t0,N3795_t1,
     N3798_t0,N3798_t1,N3801_t0,N3801_t1,N3804_t0,N3804_t1,N3834_t0,N3834_t1,N3837_t0,N3837_t1,
     N3840_t0,N3840_t1,N3843_t0,N3843_t1,N3873_t0,N3873_t1,N3876_t0,N3876_t1,N3879_t0,N3879_t1,
     N3882_t0,N3882_t1,N4193_t0,N4193_t1,N4193_t2,N4303_t0,N4303_t1,N4803_t0,N4803_t1,N4806_t0,
     N4806_t1,N4817_t0,N4817_t1,N4820_t0,N4820_t1,N4823_t0,N4823_t1,N4826_t0,N4826_t1,N4829_t0,
     N4829_t1,N4832_t0,N4832_t1,N4835_t0,N4835_t1,N4838_t0,N4838_t1,N4841_t0,N4841_t1,N4769_t0,
     N4769_t1,N4769_t2,N4769_t3,N4769_t4,N4844_t0,N4844_t1,N4847_t0,N4847_t1,N4850_t0,N4850_t1,
     N4853_t0,N4853_t1,N4856_t0,N4856_t1,N4859_t0,N4859_t1,N4862_t0,N4862_t1,N4865_t0,N4865_t1,
     N4868_t0,N4868_t1,N4874_t0,N4874_t1,N4877_t0,N4877_t1,N4880_t0,N4880_t1,N4883_t0,N4883_t1,
     N4886_t0,N4886_t1,N4889_t0,N4889_t1,N4892_t0,N4892_t1,N4895_t0,N4895_t1,N4898_t0,N4898_t1,
     N4901_t0,N4901_t1,N4904_t0,N4904_t1,N4907_t0,N4907_t1,N4910_t0,N4910_t1,N4913_t0,N4913_t1,
     N4916_t0,N4916_t1,N4919_t0,N4919_t1,N4922_t0,N4922_t1,N4925_t0,N4925_t1,N4928_t0,N4928_t1,
     N4931_t0,N4931_t1,N4934_t0,N4934_t1,N4937_t0,N4937_t1,N4940_t0,N4940_t1,N4943_t0,N4943_t1,
     N4946_t0,N4946_t1,N4949_t0,N4949_t1,N4952_t0,N4952_t1,N4955_t0,N4955_t1,N4970_t0,N4970_t1,
     N4973_t0,N4973_t1,N4976_t0,N4976_t1,N4979_t0,N4979_t1,N4982_t0,N4982_t1,N4997_t0,N4997_t1,
     N5000_t0,N5000_t1,N5003_t0,N5003_t1,N5006_t0,N5006_t1,N5009_t0,N5009_t1,N5012_t0,N5012_t1,
     N5015_t0,N5015_t1,N5018_t0,N5018_t1,N5021_t0,N5021_t1,N5024_t0,N5024_t1,N5033_t0,N5033_t1,
     N5036_t0,N5036_t1,N5039_t0,N5039_t1,N5042_t0,N5042_t1,N5049_t0,N5049_t1,N5068_t0,N5068_t1,
     N5071_t0,N5071_t1,N5074_t0,N5074_t1,N5077_t0,N5077_t1,N5080_t0,N5080_t1,N5083_t0,N5083_t1,
     N5086_t0,N5086_t1,N5089_t0,N5089_t1,N5092_t0,N5092_t1,N5095_t0,N5095_t1,N5098_t0,N5098_t1,
     N5101_t0,N5101_t1,N5104_t0,N5104_t1,N5107_t0,N5107_t1,N5114_t0,N5114_t1,N5117_t0,N5117_t1,
     N5120_t0,N5120_t1,N5123_t0,N5123_t1,N5138_t0,N5138_t1,N5141_t0,N5141_t1,N5144_t0,N5144_t1,
     N5147_t0,N5147_t1,N5150_t0,N5150_t1,N4784_t0,N4784_t1,N4790_t0,N4790_t1,N4796_t0,N4796_t1,
     N4810_t0,N4810_t1,N4814_t0,N4814_t1,N4555_t0,N4555_t1,N4555_t2,N4555_t3,N4555_t4,N4555_t5,
     N4871_t0,N4871_t1,N4586_t0,N4586_t1,N4586_t2,N4586_t3,N4586_t4,N4667_t0,N4667_t1,N4667_t2,
     N4667_t3,N4667_t4,N4667_t5,N4958_t0,N4958_t1,N4961_t0,N4961_t1,N4964_t0,N4964_t1,N4967_t0,
     N4967_t1,N4985_t0,N4985_t1,N4988_t0,N4988_t1,N4991_t0,N4991_t1,N4994_t0,N4994_t1,N5027_t0,
     N5027_t1,N4711_t0,N4711_t1,N4711_t2,N4711_t3,N4711_t4,N5030_t0,N5030_t1,N4735_t0,N4735_t1,
     N4735_t2,N4735_t3,N4735_t4,N4735_t5,N4735_t6,N5052_t0,N5052_t1,N5055_t0,N5055_t1,N5058_t0,
     N5058_t1,N5061_t0,N5061_t1,N5126_t0,N5126_t1,N5129_t0,N5129_t1,N5132_t0,N5132_t1,N5135_t0,
     N5135_t1,N5153_t0,N5153_t1,N5156_t0,N5156_t1,N5159_t0,N5159_t1,N5162_t0,N5162_t1,N5892_t0,
     N5892_t1,N5892_t2,N5892_t3,N5892_t4,N5683_t0,N5683_t1,N5683_t2,N5683_t3,N5683_t4,N5683_t5,
     N5670_t0,N5670_t1,N5670_t2,N5670_t3,N5670_t4,N5670_t5,N5670_t6,N5670_t7,N5670_t8,N5670_t9,
     N5670_t10,N5670_t11,N5654_t0,N5654_t1,N5654_t2,N5654_t3,N5654_t4,N5654_t5,N5654_t6,N5654_t7,
     N5654_t8,N5654_t9,N5654_t10,N5654_t11,N5654_t12,N5654_t13,N5654_t14,N5640_t0,N5640_t1,N5640_t2,
     N5640_t3,N5640_t4,N5640_t5,N5640_t6,N5640_t7,N5640_t8,N5640_t9,N5640_t10,N5640_t11,N5640_t12,
     N5632_t0,N5632_t1,N5632_t2,N5632_t3,N5632_t4,N5632_t5,N5632_t6,N3097_t0,N3097_t1,N3097_t2,
     N3101_t0,N3101_t1,N3101_t2,N3101_t3,N3101_t4,N3107_t0,N3107_t1,N3107_t2,N3107_t3,N3107_t4,
     N3107_t5,N5697_t0,N5697_t1,N5697_t2,N5697_t3,N5697_t4,N5697_t5,N5697_t6,N5697_t7,N5697_t8,
     N5728_t0,N5728_t1,N5728_t2,N5728_t3,N5728_t4,N5728_t5,N5707_t0,N5707_t1,N5707_t2,N5707_t3,
     N5707_t4,N5707_t5,N5707_t6,N5707_t7,N5707_t8,N5707_t9,N5690_t0,N5690_t1,N5690_t2,N5690_t3,
     N5690_t4,N5690_t5,N5718_t0,N5718_t1,N5718_t2,N5718_t3,N5718_t4,N5718_t5,N5718_t6,N5718_t7,
     N5718_t8,N3137_t0,N3137_t1,N3140_t0,N3140_t1,N3140_t2,N3144_t0,N3144_t1,N3144_t2,N3144_t3,
     N3149_t0,N3149_t1,N3149_t2,N3149_t3,N3149_t4,N5736_t0,N5736_t1,N5736_t2,N5740_t0,N5740_t1,
     N5740_t2,N5747_t0,N5747_t1,N5747_t2,N5751_t0,N5751_t1,N5751_t2,N5758_t0,N5758_t1,N5758_t2,
     N5762_t0,N5762_t1,N5762_t2,N5744_t0,N5744_t1,N5755_t0,N5755_t1,N5766_t0,N5766_t1,N5850_t0,
     N5850_t1,N5850_t2,N5850_t3,N5850_t4,N5789_t0,N5789_t1,N5789_t2,N5789_t3,N5789_t4,N5789_t5,
     N5789_t6,N5789_t7,N5789_t8,N5778_t0,N5778_t1,N5778_t2,N5778_t3,N5778_t4,N5778_t5,N5778_t6,
     N5778_t7,N5778_t8,N5778_t9,N5771_t0,N5771_t1,N5771_t2,N5771_t3,N5771_t4,N5771_t5,N3169_t0,
     N3169_t1,N3169_t2,N3173_t0,N3173_t1,N3173_t2,N3173_t3,N5856_t0,N5856_t1,N5856_t2,N5856_t3,
     N5856_t4,N5856_t5,N5837_t0,N5837_t1,N5837_t2,N5837_t3,N5837_t4,N5837_t5,N5837_t6,N5837_t7,
     N5837_t8,N5837_t9,N5837_t10,N5837_t11,N5821_t0,N5821_t1,N5821_t2,N5821_t3,N5821_t4,N5821_t5,
     N5821_t6,N5821_t7,N5821_t8,N5821_t9,N5821_t10,N5821_t11,N5821_t12,N5821_t13,N5821_t14,N5807_t0,
     N5807_t1,N5807_t2,N5807_t3,N5807_t4,N5807_t5,N5807_t6,N5807_t7,N5807_t8,N5807_t9,N5807_t10,
     N5807_t11,N5807_t12,N5799_t0,N5799_t1,N5799_t2,N5799_t3,N5799_t4,N5799_t5,N5799_t6,N3185_t0,
     N3185_t1,N3185_t2,N3189_t0,N3189_t1,N3189_t2,N3189_t3,N3189_t4,N3195_t0,N3195_t1,N3195_t2,
     N3195_t3,N3195_t4,N3195_t5,N5870_t0,N5870_t1,N5870_t2,N5870_t3,N5870_t4,N5870_t5,N5870_t6,
     N5870_t7,N5870_t8,N5870_t9,N5881_t0,N5881_t1,N5881_t2,N5881_t3,N5881_t4,N5881_t5,N5881_t6,
     N5881_t7,N5881_t8,N5881_t9,N5863_t0,N5863_t1,N5863_t2,N5863_t3,N5863_t4,N5863_t5,N3211_t0,
     N3211_t1,N3211_t2,N3215_t0,N3215_t1,N3215_t2,N3215_t3,N3215_t4,N5905_t0,N5905_t1,N5905_t2,
     N5905_t3,N5905_t4,N5905_t5,N5905_t6,N5905_t7,N5905_t8,N5936_t0,N5936_t1,N5936_t2,N5936_t3,
     N5936_t4,N5936_t5,N5915_t0,N5915_t1,N5915_t2,N5915_t3,N5915_t4,N5915_t5,N5915_t6,N5915_t7,
     N5915_t8,N5915_t9,N5898_t0,N5898_t1,N5898_t2,N5898_t3,N5898_t4,N5898_t5,N5926_t0,N5926_t1,
     N5926_t2,N5926_t3,N5926_t4,N5926_t5,N5926_t6,N5926_t7,N5926_t8,N3229_t0,N3229_t1,N3232_t0,
     N3232_t1,N3232_t2,N3236_t0,N3236_t1,N3236_t2,N3236_t3,N3241_t0,N3241_t1,N3241_t2,N3241_t3,
     N3241_t4,N6204_t0,N6204_t1,N6207_t0,N6207_t1,N6210_t0,N6210_t1,N6000_t0,N6000_t1,N5996_t0,
     N5996_t1,N5996_t2,N5991_t0,N5991_t1,N5991_t2,N5991_t3,N6018_t0,N6018_t1,N6014_t0,N6014_t1,
     N6014_t2,N6009_t0,N6009_t1,N6009_t2,N6009_t3,N6003_t0,N6003_t1,N6003_t2,N6003_t3,N6003_t4,
     N6056_t0,N6056_t1,N6052_t0,N6052_t1,N6052_t2,N6047_t0,N6047_t1,N6047_t2,N6047_t3,N6041_t0,
     N6041_t1,N6041_t2,N6041_t3,N6041_t4,N6220_t0,N6220_t1,N6079_t0,N6079_t1,N6079_t2,N6083_t0,
     N6083_t1,N6083_t2,N6087_t0,N6087_t1,N6127_t0,N6127_t1,N6127_t2,N6131_t0,N6131_t1,N6131_t2,
     N6137_t0,N6137_t1,N6137_t2,N6141_t0,N6141_t1,N6141_t2,N6145_t0,N6145_t1,N6166_t0,N6166_t1,
     N6166_t2,N6170_t0,N6170_t1,N6170_t2,N6177_t0,N6177_t1,N6177_t2,N6174_t0,N6174_t1,N6196_t0,
     N6196_t1,N6199_t0,N6199_t1,N6214_t0,N6214_t1,N6217_t0,N6217_t1,N5981_t0,N5981_t1,N5981_t2,
     N5981_t3,N5981_t4,N5981_t5,N5981_t6,N6249_t0,N6249_t1,N6252_t0,N6252_t1,N6243_t0,N6243_t1,
     N6246_t0,N6246_t1,N6232_t0,N6232_t1,N6236_t0,N6236_t1,N6263_t0,N6263_t1,N6266_t0,N6266_t1,
     N7411_t0,N7411_t1,N7414_t0,N7414_t1,N7417_t0,N7417_t1,N7420_t0,N7420_t1,N7423_t0,N7423_t1,
     N7426_t0,N7426_t1,N7429_t0,N7429_t1,N7432_t0,N7432_t1,N7435_t0,N7435_t1,N7438_t0,N7438_t1,
     N7136_t0,N7136_t1,N7136_t2,N7136_t3,N7136_t4,N6923_t0,N6923_t1,N6923_t2,N6923_t3,N6923_t4,
     N6762_t0,N6762_t1,N6762_t2,N7459_t0,N7459_t1,N7462_t0,N7462_t1,N6784_t0,N6784_t1,N6815_t0,
     N6815_t1,N6818_t0,N6818_t1,N6821_t0,N6821_t1,N6824_t0,N6824_t1,N6827_t0,N6827_t1,N6830_t0,
     N6830_t1,N6800_t0,N6800_t1,N6797_t0,N6797_t1,N6806_t0,N6806_t1,N6803_t0,N6803_t1,N6812_t0,
     N6812_t1,N6809_t0,N6809_t1,N6845_t0,N6845_t1,N7488_t0,N7488_t1,N7500_t0,N7500_t1,N7515_t0,
     N7515_t1,N7518_t0,N7518_t1,N6833_t0,N6833_t1,N6867_t0,N6867_t1,N6881_t0,N6881_t1,N7533_t0,
     N7533_t1,N7536_t0,N7536_t1,N7539_t0,N7539_t1,N7542_t0,N7542_t1,N7545_t0,N7545_t1,N7548_t0,
     N7548_t1,N6901_t0,N6901_t1,N6901_t2,N6901_t3,N6901_t4,N6901_t5,N6901_t6,N6901_t7,N6901_t8,
     N6901_t9,N6912_t0,N6912_t1,N6912_t2,N6912_t3,N6912_t4,N6912_t5,N6912_t6,N6912_t7,N6912_t8,
     N6912_t9,N6894_t0,N6894_t1,N6894_t2,N6894_t3,N6894_t4,N6894_t5,N4545_t0,N4545_t1,N4545_t2,
     N4549_t0,N4549_t1,N4549_t2,N4549_t3,N4549_t4,N6929_t0,N6929_t1,N6929_t2,N6929_t3,N6929_t4,
     N6929_t5,N4563_t0,N4563_t1,N6936_t0,N6936_t1,N6936_t2,N6936_t3,N6936_t4,N6936_t5,N6936_t6,
     N6936_t7,N6936_t8,N4566_t0,N4566_t1,N4566_t2,N6946_t0,N6946_t1,N6946_t2,N6946_t3,N6946_t4,
     N6946_t5,N6946_t6,N6946_t7,N6946_t8,N6946_t9,N4570_t0,N4570_t1,N4570_t2,N4570_t3,N6957_t0,
     N6957_t1,N6957_t2,N6957_t3,N6957_t4,N6957_t5,N6957_t6,N6957_t7,N6957_t8,N5960_t0,N5960_t1,
     N5960_t2,N5960_t3,N5960_t4,N7049_t0,N7049_t1,N7049_t2,N7049_t3,N7049_t4,N6988_t0,N6988_t1,
     N6988_t2,N6988_t3,N6988_t4,N6988_t5,N6988_t6,N6988_t7,N6988_t8,N6977_t0,N6977_t1,N6977_t2,
     N6977_t3,N6977_t4,N6977_t5,N6977_t6,N6977_t7,N6977_t8,N6977_t9,N6970_t0,N6970_t1,N6970_t2,
     N6970_t3,N6970_t4,N6970_t5,N4577_t0,N4577_t1,N4577_t2,N4581_t0,N4581_t1,N4581_t2,N4581_t3,
     N6998_t0,N6998_t1,N6998_t2,N6998_t3,N6998_t4,N6998_t5,N6998_t6,N4593_t0,N4593_t1,N4593_t2,
     N7006_t0,N7006_t1,N7006_t2,N7006_t3,N7006_t4,N7006_t5,N7006_t6,N7006_t7,N7006_t8,N7006_t9,
     N7006_t10,N7006_t11,N7006_t12,N4597_t0,N4597_t1,N4597_t2,N4597_t3,N4597_t4,N7020_t0,N7020_t1,
     N7020_t2,N7020_t3,N7020_t4,N7020_t5,N7020_t6,N7020_t7,N7020_t8,N7020_t9,N7020_t10,N7020_t11,
     N7020_t12,N7020_t13,N7020_t14,N4603_t0,N4603_t1,N4603_t2,N4603_t3,N4603_t4,N4603_t5,N7036_t0,
     N7036_t1,N7036_t2,N7036_t3,N7036_t4,N7036_t5,N7036_t6,N7036_t7,N7036_t8,N7036_t9,N7036_t10,
     N7036_t11,N7057_t0,N7057_t1,N7077_t0,N7077_t1,N7073_t0,N7073_t1,N7073_t2,N7068_t0,N7068_t1,
     N7068_t2,N7068_t3,N7095_t0,N7095_t1,N7091_t0,N7091_t1,N7091_t2,N7086_t0,N7086_t1,N7086_t2,
     N7086_t3,N7080_t0,N7080_t1,N7080_t2,N7080_t3,N7080_t4,N7100_t0,N7100_t1,N7114_t0,N7114_t1,
     N7114_t2,N7114_t3,N7114_t4,N7114_t5,N7114_t6,N7114_t7,N7114_t8,N7114_t9,N7125_t0,N7125_t1,
     N7125_t2,N7125_t3,N7125_t4,N7125_t5,N7125_t6,N7125_t7,N7125_t8,N7125_t9,N7107_t0,N7107_t1,
     N7107_t2,N7107_t3,N7107_t4,N7107_t5,N4657_t0,N4657_t1,N4657_t2,N4661_t0,N4661_t1,N4661_t2,
     N4661_t3,N4661_t4,N7149_t0,N7149_t1,N7149_t2,N7149_t3,N7149_t4,N7149_t5,N7149_t6,N7149_t7,
     N7149_t8,N7180_t0,N7180_t1,N7180_t2,N7180_t3,N7180_t4,N7180_t5,N7159_t0,N7159_t1,N7159_t2,
     N7159_t3,N7159_t4,N7159_t5,N7159_t6,N7159_t7,N7159_t8,N7159_t9,N7142_t0,N7142_t1,N7142_t2,
     N7142_t3,N7142_t4,N7142_t5,N7170_t0,N7170_t1,N7170_t2,N7170_t3,N7170_t4,N7170_t5,N7170_t6,
     N7170_t7,N7170_t8,N4675_t0,N4675_t1,N4678_t0,N4678_t1,N4678_t2,N4682_t0,N4682_t1,N4682_t2,
     N4682_t3,N4687_t0,N4687_t1,N4687_t2,N4687_t3,N4687_t4,N7194_t0,N7194_t1,N7194_t2,N7198_t0,
     N7198_t1,N7198_t2,N7205_t0,N7205_t1,N7205_t2,N7209_t0,N7209_t1,N7209_t2,N7216_t0,N7216_t1,
     N7219_t0,N7219_t1,N7202_t0,N7202_t1,N7213_t0,N7213_t1,N7191_t0,N7191_t1,N7188_t0,N7188_t1,
     N7301_t0,N7301_t1,N7301_t2,N7301_t3,N7301_t4,N7240_t0,N7240_t1,N7240_t2,N7240_t3,N7240_t4,
     N7240_t5,N7240_t6,N7240_t7,N7240_t8,N7229_t0,N7229_t1,N7229_t2,N7229_t3,N7229_t4,N7229_t5,
     N7229_t6,N7229_t7,N7229_t8,N7229_t9,N7222_t0,N7222_t1,N7222_t2,N7222_t3,N7222_t4,N7222_t5,
     N4702_t0,N4702_t1,N4702_t2,N4706_t0,N4706_t1,N4706_t2,N4706_t3,N7307_t0,N7307_t1,N7307_t2,
     N7307_t3,N7307_t4,N7307_t5,N7288_t0,N7288_t1,N7288_t2,N7288_t3,N7288_t4,N7288_t5,N7288_t6,
     N7288_t7,N7288_t8,N7288_t9,N7288_t10,N7288_t11,N7272_t0,N7272_t1,N7272_t2,N7272_t3,N7272_t4,
     N7272_t5,N7272_t6,N7272_t7,N7272_t8,N7272_t9,N7272_t10,N7272_t11,N7272_t12,N7272_t13,N7272_t14,
     N7258_t0,N7258_t1,N7258_t2,N7258_t3,N7258_t4,N7258_t5,N7258_t6,N7258_t7,N7258_t8,N7258_t9,
     N7258_t10,N7258_t11,N7258_t12,N7250_t0,N7250_t1,N7250_t2,N7250_t3,N7250_t4,N7250_t5,N7250_t6,
     N4718_t0,N4718_t1,N4718_t2,N4722_t0,N4722_t1,N4722_t2,N4722_t3,N4722_t4,N4728_t0,N4728_t1,
     N4728_t2,N4728_t3,N4728_t4,N4728_t5,N7314_t0,N7314_t1,N7314_t2,N7318_t0,N7318_t1,N7318_t2,
     N7322_t0,N7322_t1,N7331_t0,N7331_t1,N7340_t0,N7340_t1,N7343_t0,N7343_t1,N7337_t0,N7337_t1,
     N7334_t0,N7334_t1,N7355_t0,N7355_t1,N7351_t0,N7351_t1,N7351_t2,N7346_t0,N7346_t1,N7346_t2,
     N7346_t3,N7373_t0,N7373_t1,N7369_t0,N7369_t1,N7369_t2,N7364_t0,N7364_t1,N7364_t2,N7364_t3,
     N7358_t0,N7358_t1,N7358_t2,N7358_t3,N7358_t4,N7387_t0,N7387_t1,N7387_t2,N7394_t0,N7394_t1,
     N7394_t2,N7398_t0,N7398_t1,N7398_t2,N7405_t0,N7405_t1,N7408_t0,N7408_t1,N7391_t0,N7391_t1,
     N7402_t0,N7402_t1,N7381_t0,N7381_t1,N7378_t0,N7378_t1,N7441_t0,N7441_t1,N7444_t0,N7444_t1,
     N7447_t0,N7447_t1,N7450_t0,N7450_t1,N7453_t0,N7453_t1,N7456_t0,N7456_t1,N7474_t0,N7474_t1,
     N7465_t0,N7465_t1,N7468_t0,N7468_t1,N7471_t0,N7471_t1,N7479_t0,N7479_t1,N7482_t0,N7482_t1,
     N7485_t0,N7485_t1,N7491_t0,N7491_t1,N7494_t0,N7494_t1,N7497_t0,N7497_t1,N7503_t0,N7503_t1,
     N7506_t0,N7506_t1,N7509_t0,N7509_t1,N7512_t0,N7512_t1,N7530_t0,N7530_t1,N7521_t0,N7521_t1,
     N7524_t0,N7524_t1,N7527_t0,N7527_t1,N7553_t0,N7553_t1,N7574_t0,N7574_t1,N7577_t0,N7577_t1,
     N7560_t0,N7560_t1,N7563_t0,N7563_t1,N7566_t0,N7566_t1,N7569_t0,N7569_t1,N7588_t0,N7588_t1,
     N7591_t0,N7591_t1,N7582_t0,N7582_t1,N7585_t0,N7585_t1,N7620_t0,N7620_t1,N7609_t0,N7609_t1,
     N7609_t2,N7655_t0,N7655_t1,N7655_t2,N7671_t0,N7671_t1,N8196_t0,N8196_t1,N8200_t0,N8200_t1,
     N8204_t0,N8204_t1,N8208_t0,N8208_t1,N7852_t0,N7852_t1,N8114_t0,N8114_t1,N7613_t0,N7613_t1,
     N8117_t0,N8117_t1,N8131_t0,N8131_t1,N8134_t0,N8134_t1,N7650_t0,N7650_t1,N8146_t0,N8146_t1,
     N8156_t0,N8156_t1,N8166_t0,N8166_t1,N7659_t0,N7659_t1,N8169_t0,N8169_t1,N8183_t0,N8183_t1,
     N8186_t0,N8186_t1,N8580_t0,N8580_t1,N8583_t0,N8583_t1,N8586_t0,N8586_t1,N8589_t0,N8589_t1,
     N8592_t0,N8592_t1,N8595_t0,N8595_t1,N8598_t0,N8598_t1,N8601_t0,N8601_t1,N8604_t0,N8604_t1,
     N8627_t0,N8627_t1,N8333_t0,N8333_t1,N8333_t2,N8326_t0,N8326_t1,N8326_t2,N8326_t3,N8326_t4,
     N8326_t5,N8660_t0,N8660_t1,N8663_t0,N8663_t1,N8666_t0,N8666_t1,N8669_t0,N8669_t1,N8672_t0,
     N8672_t1,N8675_t0,N8675_t1,N8365_t0,N8365_t1,N8365_t2,N8358_t0,N8358_t1,N8358_t2,N8358_t3,
     N8358_t4,N8358_t5,N8687_t0,N8687_t1,N8699_t0,N8699_t1,N8711_t0,N8711_t1,N8714_t0,N8714_t1,
     N8727_t0,N8727_t1,N8730_t0,N8730_t1,N8405_t0,N8405_t1,N8405_t2,N8412_t0,N8412_t1,N8430_t0,
     N8430_t1,N8444_t0,N8444_t1,N8735_t0,N8735_t1,N8738_t0,N8738_t1,N8741_t0,N8741_t1,N8744_t0,
     N8744_t1,N8747_t0,N8747_t1,N8750_t0,N8750_t1,N8471_t0,N8471_t1,N8474_t0,N8474_t1,N8477_t0,
     N8477_t1,N8480_t0,N8480_t1,N8460_t0,N8460_t1,N8457_t0,N8457_t1,N8466_t0,N8466_t1,N8463_t0,
     N8463_t1,N8497_t0,N8497_t1,N8766_t0,N8766_t1,N8778_t0,N8778_t1,N8793_t0,N8793_t1,N8796_t0,
     N8796_t1,N8485_t0,N8485_t1,N8525_t0,N8525_t1,N8528_t0,N8528_t1,N8531_t0,N8531_t1,N8534_t0,
     N8534_t1,N8522_t0,N8522_t1,N8519_t0,N8519_t1,N7328_t0,N7328_t1,N7325_t0,N7325_t1,N8541_t0,
     N8541_t1,N8541_t2,N8548_t0,N8548_t1,N89_t0,N89_t1,N89_t2,N89_t3,N8811_t0,N8811_t1,
     N8566_t0,N8566_t1,N8569_t0,N8569_t1,N8572_t0,N8572_t1,N8575_t0,N8575_t1,N8555_t0,N8555_t1,
     N7384_t0,N7384_t1,N8561_t0,N8561_t1,N8558_t0,N8558_t1,N8678_t0,N8678_t1,N8681_t0,N8681_t1,
     N8684_t0,N8684_t1,N8690_t0,N8690_t1,N8693_t0,N8693_t1,N8696_t0,N8696_t1,N8702_t0,N8702_t1,
     N8705_t0,N8705_t1,N8708_t0,N8708_t1,N8724_t0,N8724_t1,N8718_t0,N8718_t1,N8721_t0,N8721_t1,
     N8757_t0,N8757_t1,N8760_t0,N8760_t1,N8763_t0,N8763_t1,N8769_t0,N8769_t1,N8772_t0,N8772_t1,
     N8775_t0,N8775_t1,N8781_t0,N8781_t1,N8784_t0,N8784_t1,N8787_t0,N8787_t1,N8790_t0,N8790_t1,
     N8808_t0,N8808_t1,N8799_t0,N8799_t1,N8802_t0,N8802_t1,N8805_t0,N8805_t1,N8943_t0,N8943_t1,
     N8943_t2,N8421_t0,N8421_t1,N8421_t2,N8421_t3,N8421_t4,N8421_t5,N8421_t6,N8421_t7,N8857_t0,
     N8857_t1,N8857_t2,N8871_t0,N8871_t1,N8898_t0,N8898_t1,N8898_t2,N8902_t0,N8902_t1,N9099_t0,
     N9099_t1,N9103_t0,N9103_t1,N9107_t0,N9107_t1,N9111_t0,N9111_t1,N8920_t0,N8920_t1,N8920_t2,
     N8927_t0,N8927_t1,N8927_t2,N8950_t0,N8950_t1,N8950_t2,N8956_t0,N8956_t1,N8966_t0,N8966_t1,
     N9161_t0,N9161_t1,N9165_t0,N9165_t1,N9169_t0,N9169_t1,N9173_t0,N9173_t1,N9001_t0,N9001_t1,
     N9001_t2,N9029_t0,N9029_t1,N9029_t2,N9035_t0,N9035_t1,N9068_t0,N9068_t1,N9074_t0,N9074_t1,
     N9079_t0,N9079_t1,N9083_t0,N9083_t1,N9089_t0,N9089_t1,N9095_t0,N9095_t1,N8924_t0,N8924_t1,
     N9117_t0,N9117_t1,N9127_t0,N9127_t1,N8931_t0,N8931_t1,N9146_t0,N9146_t1,N9149_t0,N9149_t1,
     N8996_t0,N8996_t1,N9183_t0,N9183_t1,N9193_t0,N9193_t1,N9203_t0,N9203_t1,N9005_t0,N9005_t1,
     N9206_t0,N9206_t1,N9220_t0,N9220_t1,N9223_t0,N9223_t1,N9268_t0,N9268_t1,N8269_t0,N8269_t1,
     N8269_t2,N8269_t3,N9408_t0,N9408_t1,N9408_t2,N9332_t0,N9332_t1,N9332_t2,N9332_t3,N9332_t4,
     N9332_t5,N8394_t0,N8394_t1,N8394_t2,N8394_t3,N8394_t4,N8394_t5,N8394_t6,N8394_t7,N8394_t8,
     N9265_t0,N9265_t1,N8262_t0,N8262_t1,N8262_t2,N8262_t3,N9423_t0,N9423_t1,N9280_t0,N9280_t1,
     N9307_t0,N9307_t1,N9307_t2,N9478_t0,N9478_t1,N9485_t0,N9485_t1,N9488_t0,N9488_t1,N9517_t0,
     N9517_t1,N9520_t0,N9520_t1,N9426_t0,N9426_t1,N9429_t0,N9429_t1,N9462_t0,N9462_t1,N9473_t0,
     N9473_t1,N9626_t0,N9626_t1,N9629_t0,N9629_t1,N9632_t0,N9632_t1,N9635_t0,N9635_t1,N9543_t0,
     N9543_t1,N9650_t0,N9650_t1,N9653_t0,N9653_t1,N9656_t0,N9656_t1,N9551_t0,N9551_t1,N9575_t0,
     N9575_t1,N9575_t2,N9698_t0,N9698_t1,N9702_t0,N9702_t1,N9608_t0,N9608_t1,N9727_t0,N9727_t1,
     N9642_t0,N9642_t1,N9646_t0,N9646_t1,N9663_t0,N9663_t1,N9667_t0,N9667_t1,N9671_t0,N9671_t1,
     N9675_t0,N9675_t1,N9679_t0,N9679_t1,N9682_t0,N9682_t1,N9685_t0,N9685_t1,N9692_t0,N9692_t1,
     N9707_t0,N9707_t1,N9711_t0,N9711_t1,N9717_t0,N9717_t1,N9723_t0,N9723_t1,N9791_t0,N9791_t1,
     N9791_t2,N8307_t0,N8307_t1,N8307_t2,N8307_t3,N8307_t4,N8307_t5,N9758_t0,N9758_t1,N9758_t2,
     N9344_t0,N9344_t1,N9344_t2,N9344_t3,N9344_t4,N9344_t5,N9754_t0,N9754_t1,N9754_t2,N9786_t0,
     N9786_t1,N9786_t2,N9820_t0,N9820_t1,N9820_t2,N9809_t0,N9809_t1,N9809_t2,N8298_t0,N8298_t1,
     N8298_t2,N8298_t3,N8298_t4,N8298_t5,N9779_t0,N9779_t1,N9779_t2,N9385_t0,N9385_t1,N9385_t2,
     N9385_t3,N9385_t4,N9385_t5,N9775_t0,N9775_t1,N9775_t2,N9817_t0,N9817_t1,N9339_t0,N9339_t1,
     N9925_t0,N9925_t1,N9925_t2,N9925_t3,N9925_t4,N9925_t5,N9932_t0,N9932_t1,N9935_t0,N9935_t1,
     N9983_t0,N9983_t1,N9986_t0,N9986_t1,N9989_t0,N9989_t1,N9992_t0,N9992_t1,N9949_t0,N9949_t1,
     N10007_t0,N10007_t1,N10010_t0,N10010_t1,N9961_t0,N9961_t1,N9964_t0,N9964_t1,N9979_t0,N9979_t1,
     N9999_t0,N9999_t1,N10003_t0,N10003_t1,N10070_t0,N10070_t1,N10073_t0,N10073_t1,N10124_t0,N10124_t1,
     N10124_t2,N10124_t3,N10124_t4,N10116_t0,N10116_t1,N10141_t0,N10141_t1,N10141_t2,N10141_t3,N10141_t4,
     N10141_t5,N10119_t0,N10119_t1,N10119_t2,N10119_t3,N10148_t0,N10148_t1,N10148_t2,N10148_t3,N10148_t4,
     N10148_t5,N10170_t0,N10170_t1,N10173_t0,N10173_t1,N10180_t0,N10180_t1,N10183_t0,N10183_t1,N10186_t0,
     N10186_t1,N10189_t0,N10189_t1,N10192_t0,N10192_t1,N10197_t0,N10197_t1,N10200_t0,N10200_t1,N10296_t0,
     N10296_t1,N10308_t0,N10308_t1,N10311_t0,N10311_t1,N10273_t0,N10273_t1,N10273_t2,N10273_t3,N10301_t0,
     N10301_t1,N10301_t2,N10301_t3,N10318_t0,N10318_t1,N10321_t0,N10321_t1,N10334_t0,N10334_t1,N10341_t0,
     N10341_t1,N10344_t0,N10344_t1,N10391_t0,N10391_t1,N10367_t0,N10367_t1,N10367_t2,N10367_t3,N10354_t0,
     N10354_t1,N10375_t0,N10375_t1,N10375_t2,N10375_t3,N10375_t4,N10406_t0,N10406_t1,N10409_t0,N10409_t1,
     N10412_t0,N10412_t1,N10415_t0,N10415_t1,N10419_t0,N10419_t1,N10422_t0,N10422_t1,N10425_t0,N10425_t1,
     N10428_t0,N10428_t1,N10399_t0,N10399_t1,N10402_t0,N10402_t1,N10388_t0,N10388_t1,N10360_t0,N10360_t1,
     N10357_t0,N10357_t1,N10381_t0,N10381_t1,N10381_t2,N10381_t3,N10381_t4,N10381_t5,N10479_t0,N10479_t1,
     N10479_t2,N10509_t0,N10509_t1,N10512_t0,N10512_t1,N10519_t0,N10519_t1,N10522_t0,N10522_t1,N10525_t0,
     N10525_t1,N10528_t0,N10528_t1,N10531_t0,N10531_t1,N10536_t0,N10536_t1,N10539_t0,N10539_t1,N10583_t0,
     N10583_t1,N10583_t2,N10589_t0,N10589_t1,N10589_t2,N10589_t3,N10602_t0,N10602_t1,N10652_t0,N10652_t1,
     N10652_t2,N10652_t3,N10652_t4,N10659_t0,N10659_t1,N10662_t0,N10662_t1,N10665_t0,N10665_t1,N10668_t0,
     N10668_t1,N10675_t0,N10675_t1,N10678_t0,N10678_t1,N10691_t0,N10691_t1,N10698_t0,N10698_t1,N10701_t0,
     N10701_t1,N10739_t0,N10739_t1,N10778_t0,N10778_t1,N10781_t0,N10781_t1,N10784_t0,N10784_t1,N10784_t2,
     N10784_t3,N10789_t0,N10789_t1,N10792_t0,N10792_t1,N10800_t0,N10800_t1,N10803_t0,N10803_t1,N10806_t0,
     N10806_t1,N10809_t0,N10809_t1,N10812_t0,N10812_t1,N10817_t0,N10817_t1,N10820_t0,N10820_t1,N10876_t0,
     N10876_t1,N10879_t0,N10879_t1,N10892_t0,N10892_t1,N10899_t0,N10899_t1,N10902_t0,N10902_t1,N10928_t0,
     N10928_t1,N10931_t0,N10931_t1,N10938_t0,N10938_t1,N10941_t0,N10941_t1,N10944_t0,N10944_t1,N10947_t0,
     N10947_t1,N10950_t0,N10950_t1,N10955_t0,N10955_t1,N10958_t0,N10958_t1,N10992_t0,N10992_t1,N10995_t0,
     N10995_t1,N11008_t0,N11008_t1,N11015_t0,N11015_t1,N11018_t0,N11018_t1,N11056_t0,N11056_t1,N11059_t0,
     N11059_t1,N11067_t0,N11067_t1,N11070_t0,N11070_t1,N11044_t0,N11044_t1,N11047_t0,N11047_t1,N11050_t0,
     N11050_t1,N11053_t0,N11053_t1,N11062_t0,N11062_t1,N11103_t0,N11103_t1,N10283_t0,N10283_t1,N10283_t2,
     N11100_t0,N11100_t1,N11124_t0,N11124_t1,N11127_t0,N11127_t1,N11130_t0,N11130_t1,N11168_t0,N11168_t1,
     N11171_t0,N11171_t1,N11174_t0,N11174_t1,N11177_t0,N11177_t1,N11159_t0,N11159_t1,N1218_t0,N1218_t1,
     N1218_t2,N11156_t0,N11156_t1,N11165_t0,N11165_t1,N10497_t0,N10497_t1,N10497_t2,N11162_t0,N11162_t1,
     N11180_t0,N11180_t1,N11205_t0,N11205_t1,N11233_t0,N11233_t1,N11236_t0,N11236_t1,N11239_t0,N11239_t1,
     N11252_t0,N11252_t1,N11257_t0,N11257_t1,N11272_t0,N11272_t1,N11302_t0,N11302_t1,N11299_t0,N11299_t1,
     N11317_t0,N11317_t1,N11323_t0,N11323_t1;
reg [3962:0] FEN;
fim PI_N53( .fault(fault), .net(N53), .FEN(FEN[0]), .op(N53_t) );
fim PI_N54( .fault(fault), .net(N54), .FEN(FEN[1]), .op(N54_t) );
fim PI_N55( .fault(fault), .net(N55), .FEN(FEN[2]), .op(N55_t) );
fim PI_N56( .fault(fault), .net(N56), .FEN(FEN[3]), .op(N56_t) );
fim PI_N57( .fault(fault), .net(N57), .FEN(FEN[4]), .op(N57_t) );
fim PI_N58( .fault(fault), .net(N58), .FEN(FEN[5]), .op(N58_t) );
fim PI_N59( .fault(fault), .net(N59), .FEN(FEN[6]), .op(N59_t) );
fim PI_N60( .fault(fault), .net(N60), .FEN(FEN[7]), .op(N60_t) );
fim PI_N61( .fault(fault), .net(N61), .FEN(FEN[8]), .op(N61_t) );
fim PI_N62( .fault(fault), .net(N62), .FEN(FEN[9]), .op(N62_t) );
fim PI_N63( .fault(fault), .net(N63), .FEN(FEN[10]), .op(N63_t) );
fim PI_N64( .fault(fault), .net(N64), .FEN(FEN[11]), .op(N64_t) );
fim PI_N65( .fault(fault), .net(N65), .FEN(FEN[12]), .op(N65_t) );
fim PI_N69( .fault(fault), .net(N69), .FEN(FEN[13]), .op(N69_t) );
fim PI_N73( .fault(fault), .net(N73), .FEN(FEN[14]), .op(N73_t) );
fim PI_N74( .fault(fault), .net(N74), .FEN(FEN[15]), .op(N74_t) );
fim PI_N75( .fault(fault), .net(N75), .FEN(FEN[16]), .op(N75_t) );
fim PI_N76( .fault(fault), .net(N76), .FEN(FEN[17]), .op(N76_t) );
fim PI_N77( .fault(fault), .net(N77), .FEN(FEN[18]), .op(N77_t) );
fim PI_N78( .fault(fault), .net(N78), .FEN(FEN[19]), .op(N78_t) );
fim PI_N79( .fault(fault), .net(N79), .FEN(FEN[20]), .op(N79_t) );
fim PI_N80( .fault(fault), .net(N80), .FEN(FEN[21]), .op(N80_t) );
fim PI_N81( .fault(fault), .net(N81), .FEN(FEN[22]), .op(N81_t) );
fim PI_N82( .fault(fault), .net(N82), .FEN(FEN[23]), .op(N82_t) );
fim PI_N83( .fault(fault), .net(N83), .FEN(FEN[24]), .op(N83_t) );
fim PI_N84( .fault(fault), .net(N84), .FEN(FEN[25]), .op(N84_t) );
fim PI_N85( .fault(fault), .net(N85), .FEN(FEN[26]), .op(N85_t) );
fim PI_N86( .fault(fault), .net(N86), .FEN(FEN[27]), .op(N86_t) );
fim PI_N87( .fault(fault), .net(N87), .FEN(FEN[28]), .op(N87_t) );
fim PI_N88( .fault(fault), .net(N88), .FEN(FEN[29]), .op(N88_t) );
fim PI_N109( .fault(fault), .net(N109), .FEN(FEN[30]), .op(N109_t) );
fim PI_N110( .fault(fault), .net(N110), .FEN(FEN[31]), .op(N110_t) );
fim PI_N111( .fault(fault), .net(N111), .FEN(FEN[32]), .op(N111_t) );
fim PI_N112( .fault(fault), .net(N112), .FEN(FEN[33]), .op(N112_t) );
fim PI_N113( .fault(fault), .net(N113), .FEN(FEN[34]), .op(N113_t) );
fim PI_N114( .fault(fault), .net(N114), .FEN(FEN[35]), .op(N114_t) );
fim PI_N133( .fault(fault), .net(N133), .FEN(FEN[36]), .op(N133_t) );
fim PI_N134( .fault(fault), .net(N134), .FEN(FEN[37]), .op(N134_t) );
fim PI_N150( .fault(fault), .net(N150), .FEN(FEN[38]), .op(N150_t) );
fim PI_N151( .fault(fault), .net(N151), .FEN(FEN[39]), .op(N151_t) );
fim PI_N152( .fault(fault), .net(N152), .FEN(FEN[40]), .op(N152_t) );
fim PI_N153( .fault(fault), .net(N153), .FEN(FEN[41]), .op(N153_t) );
fim PI_N154( .fault(fault), .net(N154), .FEN(FEN[42]), .op(N154_t) );
fim PI_N155( .fault(fault), .net(N155), .FEN(FEN[43]), .op(N155_t) );
fim PI_N156( .fault(fault), .net(N156), .FEN(FEN[44]), .op(N156_t) );
fim PI_N157( .fault(fault), .net(N157), .FEN(FEN[45]), .op(N157_t) );
fim PI_N158( .fault(fault), .net(N158), .FEN(FEN[46]), .op(N158_t) );
fim PI_N159( .fault(fault), .net(N159), .FEN(FEN[47]), .op(N159_t) );
fim PI_N160( .fault(fault), .net(N160), .FEN(FEN[48]), .op(N160_t) );
fim PI_N161( .fault(fault), .net(N161), .FEN(FEN[49]), .op(N161_t) );
fim PI_N162( .fault(fault), .net(N162), .FEN(FEN[50]), .op(N162_t) );
fim PI_N163( .fault(fault), .net(N163), .FEN(FEN[51]), .op(N163_t) );
fim PI_N164( .fault(fault), .net(N164), .FEN(FEN[52]), .op(N164_t) );
fim PI_N165( .fault(fault), .net(N165), .FEN(FEN[53]), .op(N165_t) );
fim PI_N166( .fault(fault), .net(N166), .FEN(FEN[54]), .op(N166_t) );
fim PI_N167( .fault(fault), .net(N167), .FEN(FEN[55]), .op(N167_t) );
fim PI_N168( .fault(fault), .net(N168), .FEN(FEN[56]), .op(N168_t) );
fim PI_N169( .fault(fault), .net(N169), .FEN(FEN[57]), .op(N169_t) );
fim PI_N170( .fault(fault), .net(N170), .FEN(FEN[58]), .op(N170_t) );
fim PI_N171( .fault(fault), .net(N171), .FEN(FEN[59]), .op(N171_t) );
fim PI_N172( .fault(fault), .net(N172), .FEN(FEN[60]), .op(N172_t) );
fim PI_N173( .fault(fault), .net(N173), .FEN(FEN[61]), .op(N173_t) );
fim PI_N174( .fault(fault), .net(N174), .FEN(FEN[62]), .op(N174_t) );
fim PI_N175( .fault(fault), .net(N175), .FEN(FEN[63]), .op(N175_t) );
fim PI_N176( .fault(fault), .net(N176), .FEN(FEN[64]), .op(N176_t) );
fim PI_N177( .fault(fault), .net(N177), .FEN(FEN[65]), .op(N177_t) );
fim PI_N178( .fault(fault), .net(N178), .FEN(FEN[66]), .op(N178_t) );
fim PI_N179( .fault(fault), .net(N179), .FEN(FEN[67]), .op(N179_t) );
fim PI_N180( .fault(fault), .net(N180), .FEN(FEN[68]), .op(N180_t) );
fim PI_N181( .fault(fault), .net(N181), .FEN(FEN[69]), .op(N181_t) );
fim PI_N182( .fault(fault), .net(N182), .FEN(FEN[70]), .op(N182_t) );
fim PI_N183( .fault(fault), .net(N183), .FEN(FEN[71]), .op(N183_t) );
fim PI_N184( .fault(fault), .net(N184), .FEN(FEN[72]), .op(N184_t) );
fim PI_N185( .fault(fault), .net(N185), .FEN(FEN[73]), .op(N185_t) );
fim PI_N186( .fault(fault), .net(N186), .FEN(FEN[74]), .op(N186_t) );
fim PI_N187( .fault(fault), .net(N187), .FEN(FEN[75]), .op(N187_t) );
fim PI_N188( .fault(fault), .net(N188), .FEN(FEN[76]), .op(N188_t) );
fim PI_N189( .fault(fault), .net(N189), .FEN(FEN[77]), .op(N189_t) );
fim PI_N190( .fault(fault), .net(N190), .FEN(FEN[78]), .op(N190_t) );
fim PI_N191( .fault(fault), .net(N191), .FEN(FEN[79]), .op(N191_t) );
fim PI_N192( .fault(fault), .net(N192), .FEN(FEN[80]), .op(N192_t) );
fim PI_N193( .fault(fault), .net(N193), .FEN(FEN[81]), .op(N193_t) );
fim PI_N194( .fault(fault), .net(N194), .FEN(FEN[82]), .op(N194_t) );
fim PI_N195( .fault(fault), .net(N195), .FEN(FEN[83]), .op(N195_t) );
fim PI_N196( .fault(fault), .net(N196), .FEN(FEN[84]), .op(N196_t) );
fim PI_N197( .fault(fault), .net(N197), .FEN(FEN[85]), .op(N197_t) );
fim PI_N198( .fault(fault), .net(N198), .FEN(FEN[86]), .op(N198_t) );
fim PI_N199( .fault(fault), .net(N199), .FEN(FEN[87]), .op(N199_t) );
fim PI_N200( .fault(fault), .net(N200), .FEN(FEN[88]), .op(N200_t) );
fim PI_N201( .fault(fault), .net(N201), .FEN(FEN[89]), .op(N201_t) );
fim PI_N202( .fault(fault), .net(N202), .FEN(FEN[90]), .op(N202_t) );
fim PI_N203( .fault(fault), .net(N203), .FEN(FEN[91]), .op(N203_t) );
fim PI_N204( .fault(fault), .net(N204), .FEN(FEN[92]), .op(N204_t) );
fim PI_N205( .fault(fault), .net(N205), .FEN(FEN[93]), .op(N205_t) );
fim PI_N206( .fault(fault), .net(N206), .FEN(FEN[94]), .op(N206_t) );
fim PI_N207( .fault(fault), .net(N207), .FEN(FEN[95]), .op(N207_t) );
fim PI_N208( .fault(fault), .net(N208), .FEN(FEN[96]), .op(N208_t) );
fim PI_N209( .fault(fault), .net(N209), .FEN(FEN[97]), .op(N209_t) );
fim PI_N210( .fault(fault), .net(N210), .FEN(FEN[98]), .op(N210_t) );
fim PI_N211( .fault(fault), .net(N211), .FEN(FEN[99]), .op(N211_t) );
fim PI_N212( .fault(fault), .net(N212), .FEN(FEN[100]), .op(N212_t) );
fim PI_N213( .fault(fault), .net(N213), .FEN(FEN[101]), .op(N213_t) );
fim PI_N214( .fault(fault), .net(N214), .FEN(FEN[102]), .op(N214_t) );
fim PI_N215( .fault(fault), .net(N215), .FEN(FEN[103]), .op(N215_t) );
fim PI_N216( .fault(fault), .net(N216), .FEN(FEN[104]), .op(N216_t) );
fim PI_N217( .fault(fault), .net(N217), .FEN(FEN[105]), .op(N217_t) );
fim PI_N218( .fault(fault), .net(N218), .FEN(FEN[106]), .op(N218_t) );
fim PI_N219( .fault(fault), .net(N219), .FEN(FEN[107]), .op(N219_t) );
fim PI_N220( .fault(fault), .net(N220), .FEN(FEN[108]), .op(N220_t) );
fim PI_N221( .fault(fault), .net(N221), .FEN(FEN[109]), .op(N221_t) );
fim PI_N222( .fault(fault), .net(N222), .FEN(FEN[110]), .op(N222_t) );
fim PI_N223( .fault(fault), .net(N223), .FEN(FEN[111]), .op(N223_t) );
fim PI_N224( .fault(fault), .net(N224), .FEN(FEN[112]), .op(N224_t) );
fim PI_N225( .fault(fault), .net(N225), .FEN(FEN[113]), .op(N225_t) );
fim PI_N226( .fault(fault), .net(N226), .FEN(FEN[114]), .op(N226_t) );
fim PI_N227( .fault(fault), .net(N227), .FEN(FEN[115]), .op(N227_t) );
fim PI_N228( .fault(fault), .net(N228), .FEN(FEN[116]), .op(N228_t) );
fim PI_N229( .fault(fault), .net(N229), .FEN(FEN[117]), .op(N229_t) );
fim PI_N230( .fault(fault), .net(N230), .FEN(FEN[118]), .op(N230_t) );
fim PI_N231( .fault(fault), .net(N231), .FEN(FEN[119]), .op(N231_t) );
fim PI_N232( .fault(fault), .net(N232), .FEN(FEN[120]), .op(N232_t) );
fim PI_N233( .fault(fault), .net(N233), .FEN(FEN[121]), .op(N233_t) );
fim PI_N234( .fault(fault), .net(N234), .FEN(FEN[122]), .op(N234_t) );
fim PI_N235( .fault(fault), .net(N235), .FEN(FEN[123]), .op(N235_t) );
fim PI_N236( .fault(fault), .net(N236), .FEN(FEN[124]), .op(N236_t) );
fim PI_N237( .fault(fault), .net(N237), .FEN(FEN[125]), .op(N237_t) );
fim PI_N238( .fault(fault), .net(N238), .FEN(FEN[126]), .op(N238_t) );
fim PI_N239( .fault(fault), .net(N239), .FEN(FEN[127]), .op(N239_t) );
fim PI_N240( .fault(fault), .net(N240), .FEN(FEN[128]), .op(N240_t) );
fim PI_N241_I( .fault(fault), .net(N241_I), .FEN(FEN[129]), .op(N241_I_t) );
fim FAN_N1_0 ( .fault(fault), .net(N1), .FEN(FEN[130]), .op(N1_t0) );
fim FAN_N1_1 ( .fault(fault), .net(N1), .FEN(FEN[131]), .op(N1_t1) );
fim FAN_N1_2 ( .fault(fault), .net(N1), .FEN(FEN[132]), .op(N1_t2) );
fim FAN_N248_0 ( .fault(fault), .net(N248), .FEN(FEN[133]), .op(N248_t0) );
fim FAN_N248_1 ( .fault(fault), .net(N248), .FEN(FEN[134]), .op(N248_t1) );
fim FAN_N254_0 ( .fault(fault), .net(N254), .FEN(FEN[135]), .op(N254_t0) );
fim FAN_N254_1 ( .fault(fault), .net(N254), .FEN(FEN[136]), .op(N254_t1) );
fim FAN_N257_0 ( .fault(fault), .net(N257), .FEN(FEN[137]), .op(N257_t0) );
fim FAN_N257_1 ( .fault(fault), .net(N257), .FEN(FEN[138]), .op(N257_t1) );
fim FAN_N260_0 ( .fault(fault), .net(N260), .FEN(FEN[139]), .op(N260_t0) );
fim FAN_N260_1 ( .fault(fault), .net(N260), .FEN(FEN[140]), .op(N260_t1) );
fim FAN_N263_0 ( .fault(fault), .net(N263), .FEN(FEN[141]), .op(N263_t0) );
fim FAN_N263_1 ( .fault(fault), .net(N263), .FEN(FEN[142]), .op(N263_t1) );
fim FAN_N263_2 ( .fault(fault), .net(N263), .FEN(FEN[143]), .op(N263_t2) );
fim FAN_N267_0 ( .fault(fault), .net(N267), .FEN(FEN[144]), .op(N267_t0) );
fim FAN_N267_1 ( .fault(fault), .net(N267), .FEN(FEN[145]), .op(N267_t1) );
fim FAN_N267_2 ( .fault(fault), .net(N267), .FEN(FEN[146]), .op(N267_t2) );
fim FAN_N274_0 ( .fault(fault), .net(N274), .FEN(FEN[147]), .op(N274_t0) );
fim FAN_N274_1 ( .fault(fault), .net(N274), .FEN(FEN[148]), .op(N274_t1) );
fim FAN_N280_0 ( .fault(fault), .net(N280), .FEN(FEN[149]), .op(N280_t0) );
fim FAN_N280_1 ( .fault(fault), .net(N280), .FEN(FEN[150]), .op(N280_t1) );
fim FAN_N283_0 ( .fault(fault), .net(N283), .FEN(FEN[151]), .op(N283_t0) );
fim FAN_N283_1 ( .fault(fault), .net(N283), .FEN(FEN[152]), .op(N283_t1) );
fim FAN_N286_0 ( .fault(fault), .net(N286), .FEN(FEN[153]), .op(N286_t0) );
fim FAN_N286_1 ( .fault(fault), .net(N286), .FEN(FEN[154]), .op(N286_t1) );
fim FAN_N289_0 ( .fault(fault), .net(N289), .FEN(FEN[155]), .op(N289_t0) );
fim FAN_N289_1 ( .fault(fault), .net(N289), .FEN(FEN[156]), .op(N289_t1) );
fim FAN_N289_2 ( .fault(fault), .net(N289), .FEN(FEN[157]), .op(N289_t2) );
fim FAN_N293_0 ( .fault(fault), .net(N293), .FEN(FEN[158]), .op(N293_t0) );
fim FAN_N293_1 ( .fault(fault), .net(N293), .FEN(FEN[159]), .op(N293_t1) );
fim FAN_N296_0 ( .fault(fault), .net(N296), .FEN(FEN[160]), .op(N296_t0) );
fim FAN_N296_1 ( .fault(fault), .net(N296), .FEN(FEN[161]), .op(N296_t1) );
fim FAN_N299_0 ( .fault(fault), .net(N299), .FEN(FEN[162]), .op(N299_t0) );
fim FAN_N299_1 ( .fault(fault), .net(N299), .FEN(FEN[163]), .op(N299_t1) );
fim FAN_N299_2 ( .fault(fault), .net(N299), .FEN(FEN[164]), .op(N299_t2) );
fim FAN_N303_0 ( .fault(fault), .net(N303), .FEN(FEN[165]), .op(N303_t0) );
fim FAN_N303_1 ( .fault(fault), .net(N303), .FEN(FEN[166]), .op(N303_t1) );
fim FAN_N303_2 ( .fault(fault), .net(N303), .FEN(FEN[167]), .op(N303_t2) );
fim FAN_N307_0 ( .fault(fault), .net(N307), .FEN(FEN[168]), .op(N307_t0) );
fim FAN_N307_1 ( .fault(fault), .net(N307), .FEN(FEN[169]), .op(N307_t1) );
fim FAN_N310_0 ( .fault(fault), .net(N310), .FEN(FEN[170]), .op(N310_t0) );
fim FAN_N310_1 ( .fault(fault), .net(N310), .FEN(FEN[171]), .op(N310_t1) );
fim FAN_N313_0 ( .fault(fault), .net(N313), .FEN(FEN[172]), .op(N313_t0) );
fim FAN_N313_1 ( .fault(fault), .net(N313), .FEN(FEN[173]), .op(N313_t1) );
fim FAN_N316_0 ( .fault(fault), .net(N316), .FEN(FEN[174]), .op(N316_t0) );
fim FAN_N316_1 ( .fault(fault), .net(N316), .FEN(FEN[175]), .op(N316_t1) );
fim FAN_N319_0 ( .fault(fault), .net(N319), .FEN(FEN[176]), .op(N319_t0) );
fim FAN_N319_1 ( .fault(fault), .net(N319), .FEN(FEN[177]), .op(N319_t1) );
fim FAN_N322_0 ( .fault(fault), .net(N322), .FEN(FEN[178]), .op(N322_t0) );
fim FAN_N322_1 ( .fault(fault), .net(N322), .FEN(FEN[179]), .op(N322_t1) );
fim FAN_N325_0 ( .fault(fault), .net(N325), .FEN(FEN[180]), .op(N325_t0) );
fim FAN_N325_1 ( .fault(fault), .net(N325), .FEN(FEN[181]), .op(N325_t1) );
fim FAN_N328_0 ( .fault(fault), .net(N328), .FEN(FEN[182]), .op(N328_t0) );
fim FAN_N328_1 ( .fault(fault), .net(N328), .FEN(FEN[183]), .op(N328_t1) );
fim FAN_N331_0 ( .fault(fault), .net(N331), .FEN(FEN[184]), .op(N331_t0) );
fim FAN_N331_1 ( .fault(fault), .net(N331), .FEN(FEN[185]), .op(N331_t1) );
fim FAN_N334_0 ( .fault(fault), .net(N334), .FEN(FEN[186]), .op(N334_t0) );
fim FAN_N334_1 ( .fault(fault), .net(N334), .FEN(FEN[187]), .op(N334_t1) );
fim FAN_N337_0 ( .fault(fault), .net(N337), .FEN(FEN[188]), .op(N337_t0) );
fim FAN_N337_1 ( .fault(fault), .net(N337), .FEN(FEN[189]), .op(N337_t1) );
fim FAN_N343_0 ( .fault(fault), .net(N343), .FEN(FEN[190]), .op(N343_t0) );
fim FAN_N343_1 ( .fault(fault), .net(N343), .FEN(FEN[191]), .op(N343_t1) );
fim FAN_N346_0 ( .fault(fault), .net(N346), .FEN(FEN[192]), .op(N346_t0) );
fim FAN_N346_1 ( .fault(fault), .net(N346), .FEN(FEN[193]), .op(N346_t1) );
fim FAN_N349_0 ( .fault(fault), .net(N349), .FEN(FEN[194]), .op(N349_t0) );
fim FAN_N349_1 ( .fault(fault), .net(N349), .FEN(FEN[195]), .op(N349_t1) );
fim FAN_N352_0 ( .fault(fault), .net(N352), .FEN(FEN[196]), .op(N352_t0) );
fim FAN_N352_1 ( .fault(fault), .net(N352), .FEN(FEN[197]), .op(N352_t1) );
fim FAN_N355_0 ( .fault(fault), .net(N355), .FEN(FEN[198]), .op(N355_t0) );
fim FAN_N355_1 ( .fault(fault), .net(N355), .FEN(FEN[199]), .op(N355_t1) );
fim FAN_N358_0 ( .fault(fault), .net(N358), .FEN(FEN[200]), .op(N358_t0) );
fim FAN_N358_1 ( .fault(fault), .net(N358), .FEN(FEN[201]), .op(N358_t1) );
fim FAN_N361_0 ( .fault(fault), .net(N361), .FEN(FEN[202]), .op(N361_t0) );
fim FAN_N361_1 ( .fault(fault), .net(N361), .FEN(FEN[203]), .op(N361_t1) );
fim FAN_N364_0 ( .fault(fault), .net(N364), .FEN(FEN[204]), .op(N364_t0) );
fim FAN_N364_1 ( .fault(fault), .net(N364), .FEN(FEN[205]), .op(N364_t1) );
fim FAN_N15_0 ( .fault(fault), .net(N15), .FEN(FEN[206]), .op(N15_t0) );
fim FAN_N15_1 ( .fault(fault), .net(N15), .FEN(FEN[207]), .op(N15_t1) );
fim FAN_N5_0 ( .fault(fault), .net(N5), .FEN(FEN[208]), .op(N5_t0) );
fim FAN_N5_1 ( .fault(fault), .net(N5), .FEN(FEN[209]), .op(N5_t1) );
fim FAN_N5_2 ( .fault(fault), .net(N5), .FEN(FEN[210]), .op(N5_t2) );
fim FAN_N38_0 ( .fault(fault), .net(N38), .FEN(FEN[211]), .op(N38_t0) );
fim FAN_N38_1 ( .fault(fault), .net(N38), .FEN(FEN[212]), .op(N38_t1) );
fim FAN_N12_0 ( .fault(fault), .net(N12), .FEN(FEN[213]), .op(N12_t0) );
fim FAN_N12_1 ( .fault(fault), .net(N12), .FEN(FEN[214]), .op(N12_t1) );
fim FAN_N9_0 ( .fault(fault), .net(N9), .FEN(FEN[215]), .op(N9_t0) );
fim FAN_N9_1 ( .fault(fault), .net(N9), .FEN(FEN[216]), .op(N9_t1) );
fim FAN_N245_0 ( .fault(fault), .net(N245), .FEN(FEN[217]), .op(N245_t0) );
fim FAN_N245_1 ( .fault(fault), .net(N245), .FEN(FEN[218]), .op(N245_t1) );
fim FAN_N251_0 ( .fault(fault), .net(N251), .FEN(FEN[219]), .op(N251_t0) );
fim FAN_N251_1 ( .fault(fault), .net(N251), .FEN(FEN[220]), .op(N251_t1) );
fim FAN_N106_0 ( .fault(fault), .net(N106), .FEN(FEN[221]), .op(N106_t0) );
fim FAN_N106_1 ( .fault(fault), .net(N106), .FEN(FEN[222]), .op(N106_t1) );
fim FAN_N18_0 ( .fault(fault), .net(N18), .FEN(FEN[223]), .op(N18_t0) );
fim FAN_N18_1 ( .fault(fault), .net(N18), .FEN(FEN[224]), .op(N18_t1) );
fim FAN_N18_2 ( .fault(fault), .net(N18), .FEN(FEN[225]), .op(N18_t2) );
fim FAN_N18_3 ( .fault(fault), .net(N18), .FEN(FEN[226]), .op(N18_t3) );
fim FAN_N382_0 ( .fault(fault), .net(N382), .FEN(FEN[227]), .op(N382_t0) );
fim FAN_N382_1 ( .fault(fault), .net(N382), .FEN(FEN[228]), .op(N382_t1) );
fim FAN_N382_2 ( .fault(fault), .net(N382), .FEN(FEN[229]), .op(N382_t2) );
fim FAN_N382_3 ( .fault(fault), .net(N382), .FEN(FEN[230]), .op(N382_t3) );
fim FAN_N271_0 ( .fault(fault), .net(N271), .FEN(FEN[231]), .op(N271_t0) );
fim FAN_N271_1 ( .fault(fault), .net(N271), .FEN(FEN[232]), .op(N271_t1) );
fim FAN_N277_0 ( .fault(fault), .net(N277), .FEN(FEN[233]), .op(N277_t0) );
fim FAN_N277_1 ( .fault(fault), .net(N277), .FEN(FEN[234]), .op(N277_t1) );
fim FAN_N367_0 ( .fault(fault), .net(N367), .FEN(FEN[235]), .op(N367_t0) );
fim FAN_N367_1 ( .fault(fault), .net(N367), .FEN(FEN[236]), .op(N367_t1) );
fim FAN_N367_2 ( .fault(fault), .net(N367), .FEN(FEN[237]), .op(N367_t2) );
fim FAN_N367_3 ( .fault(fault), .net(N367), .FEN(FEN[238]), .op(N367_t3) );
fim FAN_N367_4 ( .fault(fault), .net(N367), .FEN(FEN[239]), .op(N367_t4) );
fim FAN_N367_5 ( .fault(fault), .net(N367), .FEN(FEN[240]), .op(N367_t5) );
fim FAN_N367_6 ( .fault(fault), .net(N367), .FEN(FEN[241]), .op(N367_t6) );
fim FAN_N367_7 ( .fault(fault), .net(N367), .FEN(FEN[242]), .op(N367_t7) );
fim FAN_N367_8 ( .fault(fault), .net(N367), .FEN(FEN[243]), .op(N367_t8) );
fim FAN_N367_9 ( .fault(fault), .net(N367), .FEN(FEN[244]), .op(N367_t9) );
fim FAN_N367_10 ( .fault(fault), .net(N367), .FEN(FEN[245]), .op(N367_t10) );
fim FAN_N367_11 ( .fault(fault), .net(N367), .FEN(FEN[246]), .op(N367_t11) );
fim FAN_N367_12 ( .fault(fault), .net(N367), .FEN(FEN[247]), .op(N367_t12) );
fim FAN_N367_13 ( .fault(fault), .net(N367), .FEN(FEN[248]), .op(N367_t13) );
fim FAN_N340_0 ( .fault(fault), .net(N340), .FEN(FEN[249]), .op(N340_t0) );
fim FAN_N340_1 ( .fault(fault), .net(N340), .FEN(FEN[250]), .op(N340_t1) );
fim FAN_N528_0 ( .fault(fault), .net(N528), .FEN(FEN[251]), .op(N528_t0) );
fim FAN_N528_1 ( .fault(fault), .net(N528), .FEN(FEN[252]), .op(N528_t1) );
fim FAN_N578_0 ( .fault(fault), .net(N578), .FEN(FEN[253]), .op(N578_t0) );
fim FAN_N578_1 ( .fault(fault), .net(N578), .FEN(FEN[254]), .op(N578_t1) );
fim FAN_N575_0 ( .fault(fault), .net(N575), .FEN(FEN[255]), .op(N575_t0) );
fim FAN_N575_1 ( .fault(fault), .net(N575), .FEN(FEN[256]), .op(N575_t1) );
fim FAN_N494_0 ( .fault(fault), .net(N494), .FEN(FEN[257]), .op(N494_t0) );
fim FAN_N494_1 ( .fault(fault), .net(N494), .FEN(FEN[258]), .op(N494_t1) );
fim FAN_N590_0 ( .fault(fault), .net(N590), .FEN(FEN[259]), .op(N590_t0) );
fim FAN_N590_1 ( .fault(fault), .net(N590), .FEN(FEN[260]), .op(N590_t1) );
fim FAN_N657_0 ( .fault(fault), .net(N657), .FEN(FEN[261]), .op(N657_t0) );
fim FAN_N657_1 ( .fault(fault), .net(N657), .FEN(FEN[262]), .op(N657_t1) );
fim FAN_N469_0 ( .fault(fault), .net(N469), .FEN(FEN[263]), .op(N469_t0) );
fim FAN_N469_1 ( .fault(fault), .net(N469), .FEN(FEN[264]), .op(N469_t1) );
fim FAN_N596_0 ( .fault(fault), .net(N596), .FEN(FEN[265]), .op(N596_t0) );
fim FAN_N596_1 ( .fault(fault), .net(N596), .FEN(FEN[266]), .op(N596_t1) );
fim FAN_N242_0 ( .fault(fault), .net(N242), .FEN(FEN[267]), .op(N242_t0) );
fim FAN_N242_1 ( .fault(fault), .net(N242), .FEN(FEN[268]), .op(N242_t1) );
fim FAN_N593_0 ( .fault(fault), .net(N593), .FEN(FEN[269]), .op(N593_t0) );
fim FAN_N593_1 ( .fault(fault), .net(N593), .FEN(FEN[270]), .op(N593_t1) );
fim FAN_N625_0 ( .fault(fault), .net(N625), .FEN(FEN[271]), .op(N625_t0) );
fim FAN_N625_1 ( .fault(fault), .net(N625), .FEN(FEN[272]), .op(N625_t1) );
fim FAN_N871_0 ( .fault(fault), .net(N871), .FEN(FEN[273]), .op(N871_t0) );
fim FAN_N871_1 ( .fault(fault), .net(N871), .FEN(FEN[274]), .op(N871_t1) );
fim FAN_N628_0 ( .fault(fault), .net(N628), .FEN(FEN[275]), .op(N628_t0) );
fim FAN_N628_1 ( .fault(fault), .net(N628), .FEN(FEN[276]), .op(N628_t1) );
fim FAN_N628_2 ( .fault(fault), .net(N628), .FEN(FEN[277]), .op(N628_t2) );
fim FAN_N682_0 ( .fault(fault), .net(N682), .FEN(FEN[278]), .op(N682_t0) );
fim FAN_N682_1 ( .fault(fault), .net(N682), .FEN(FEN[279]), .op(N682_t1) );
fim FAN_N682_2 ( .fault(fault), .net(N682), .FEN(FEN[280]), .op(N682_t2) );
fim FAN_N682_3 ( .fault(fault), .net(N682), .FEN(FEN[281]), .op(N682_t3) );
fim FAN_N682_4 ( .fault(fault), .net(N682), .FEN(FEN[282]), .op(N682_t4) );
fim FAN_N632_0 ( .fault(fault), .net(N632), .FEN(FEN[283]), .op(N632_t0) );
fim FAN_N632_1 ( .fault(fault), .net(N632), .FEN(FEN[284]), .op(N632_t1) );
fim FAN_N632_2 ( .fault(fault), .net(N632), .FEN(FEN[285]), .op(N632_t2) );
fim FAN_N676_0 ( .fault(fault), .net(N676), .FEN(FEN[286]), .op(N676_t0) );
fim FAN_N676_1 ( .fault(fault), .net(N676), .FEN(FEN[287]), .op(N676_t1) );
fim FAN_N676_2 ( .fault(fault), .net(N676), .FEN(FEN[288]), .op(N676_t2) );
fim FAN_N676_3 ( .fault(fault), .net(N676), .FEN(FEN[289]), .op(N676_t3) );
fim FAN_N676_4 ( .fault(fault), .net(N676), .FEN(FEN[290]), .op(N676_t4) );
fim FAN_N700_0 ( .fault(fault), .net(N700), .FEN(FEN[291]), .op(N700_t0) );
fim FAN_N700_1 ( .fault(fault), .net(N700), .FEN(FEN[292]), .op(N700_t1) );
fim FAN_N700_2 ( .fault(fault), .net(N700), .FEN(FEN[293]), .op(N700_t2) );
fim FAN_N700_3 ( .fault(fault), .net(N700), .FEN(FEN[294]), .op(N700_t3) );
fim FAN_N614_0 ( .fault(fault), .net(N614), .FEN(FEN[295]), .op(N614_t0) );
fim FAN_N614_1 ( .fault(fault), .net(N614), .FEN(FEN[296]), .op(N614_t1) );
fim FAN_N614_2 ( .fault(fault), .net(N614), .FEN(FEN[297]), .op(N614_t2) );
fim FAN_N614_3 ( .fault(fault), .net(N614), .FEN(FEN[298]), .op(N614_t3) );
fim FAN_N614_4 ( .fault(fault), .net(N614), .FEN(FEN[299]), .op(N614_t4) );
fim FAN_N614_5 ( .fault(fault), .net(N614), .FEN(FEN[300]), .op(N614_t5) );
fim FAN_N614_6 ( .fault(fault), .net(N614), .FEN(FEN[301]), .op(N614_t6) );
fim FAN_N614_7 ( .fault(fault), .net(N614), .FEN(FEN[302]), .op(N614_t7) );
fim FAN_N614_8 ( .fault(fault), .net(N614), .FEN(FEN[303]), .op(N614_t8) );
fim FAN_N614_9 ( .fault(fault), .net(N614), .FEN(FEN[304]), .op(N614_t9) );
fim FAN_N689_0 ( .fault(fault), .net(N689), .FEN(FEN[305]), .op(N689_t0) );
fim FAN_N689_1 ( .fault(fault), .net(N689), .FEN(FEN[306]), .op(N689_t1) );
fim FAN_N689_2 ( .fault(fault), .net(N689), .FEN(FEN[307]), .op(N689_t2) );
fim FAN_N689_3 ( .fault(fault), .net(N689), .FEN(FEN[308]), .op(N689_t3) );
fim FAN_N689_4 ( .fault(fault), .net(N689), .FEN(FEN[309]), .op(N689_t4) );
fim FAN_N695_0 ( .fault(fault), .net(N695), .FEN(FEN[310]), .op(N695_t0) );
fim FAN_N695_1 ( .fault(fault), .net(N695), .FEN(FEN[311]), .op(N695_t1) );
fim FAN_N695_2 ( .fault(fault), .net(N695), .FEN(FEN[312]), .op(N695_t2) );
fim FAN_N695_3 ( .fault(fault), .net(N695), .FEN(FEN[313]), .op(N695_t3) );
fim FAN_N750_0 ( .fault(fault), .net(N750), .FEN(FEN[314]), .op(N750_t0) );
fim FAN_N750_1 ( .fault(fault), .net(N750), .FEN(FEN[315]), .op(N750_t1) );
fim FAN_N750_2 ( .fault(fault), .net(N750), .FEN(FEN[316]), .op(N750_t2) );
fim FAN_N750_3 ( .fault(fault), .net(N750), .FEN(FEN[317]), .op(N750_t3) );
fim FAN_N666_0 ( .fault(fault), .net(N666), .FEN(FEN[318]), .op(N666_t0) );
fim FAN_N666_1 ( .fault(fault), .net(N666), .FEN(FEN[319]), .op(N666_t1) );
fim FAN_N666_2 ( .fault(fault), .net(N666), .FEN(FEN[320]), .op(N666_t2) );
fim FAN_N666_3 ( .fault(fault), .net(N666), .FEN(FEN[321]), .op(N666_t3) );
fim FAN_N666_4 ( .fault(fault), .net(N666), .FEN(FEN[322]), .op(N666_t4) );
fim FAN_N660_0 ( .fault(fault), .net(N660), .FEN(FEN[323]), .op(N660_t0) );
fim FAN_N660_1 ( .fault(fault), .net(N660), .FEN(FEN[324]), .op(N660_t1) );
fim FAN_N660_2 ( .fault(fault), .net(N660), .FEN(FEN[325]), .op(N660_t2) );
fim FAN_N660_3 ( .fault(fault), .net(N660), .FEN(FEN[326]), .op(N660_t3) );
fim FAN_N660_4 ( .fault(fault), .net(N660), .FEN(FEN[327]), .op(N660_t4) );
fim FAN_N651_0 ( .fault(fault), .net(N651), .FEN(FEN[328]), .op(N651_t0) );
fim FAN_N651_1 ( .fault(fault), .net(N651), .FEN(FEN[329]), .op(N651_t1) );
fim FAN_N651_2 ( .fault(fault), .net(N651), .FEN(FEN[330]), .op(N651_t2) );
fim FAN_N651_3 ( .fault(fault), .net(N651), .FEN(FEN[331]), .op(N651_t3) );
fim FAN_N651_4 ( .fault(fault), .net(N651), .FEN(FEN[332]), .op(N651_t4) );
fim FAN_N644_0 ( .fault(fault), .net(N644), .FEN(FEN[333]), .op(N644_t0) );
fim FAN_N644_1 ( .fault(fault), .net(N644), .FEN(FEN[334]), .op(N644_t1) );
fim FAN_N644_2 ( .fault(fault), .net(N644), .FEN(FEN[335]), .op(N644_t2) );
fim FAN_N644_3 ( .fault(fault), .net(N644), .FEN(FEN[336]), .op(N644_t3) );
fim FAN_N644_4 ( .fault(fault), .net(N644), .FEN(FEN[337]), .op(N644_t4) );
fim FAN_N644_5 ( .fault(fault), .net(N644), .FEN(FEN[338]), .op(N644_t5) );
fim FAN_N609_0 ( .fault(fault), .net(N609), .FEN(FEN[339]), .op(N609_t0) );
fim FAN_N609_1 ( .fault(fault), .net(N609), .FEN(FEN[340]), .op(N609_t1) );
fim FAN_N609_2 ( .fault(fault), .net(N609), .FEN(FEN[341]), .op(N609_t2) );
fim FAN_N609_3 ( .fault(fault), .net(N609), .FEN(FEN[342]), .op(N609_t3) );
fim FAN_N604_0 ( .fault(fault), .net(N604), .FEN(FEN[343]), .op(N604_t0) );
fim FAN_N604_1 ( .fault(fault), .net(N604), .FEN(FEN[344]), .op(N604_t1) );
fim FAN_N604_2 ( .fault(fault), .net(N604), .FEN(FEN[345]), .op(N604_t2) );
fim FAN_N604_3 ( .fault(fault), .net(N604), .FEN(FEN[346]), .op(N604_t3) );
fim FAN_N742_0 ( .fault(fault), .net(N742), .FEN(FEN[347]), .op(N742_t0) );
fim FAN_N742_1 ( .fault(fault), .net(N742), .FEN(FEN[348]), .op(N742_t1) );
fim FAN_N742_2 ( .fault(fault), .net(N742), .FEN(FEN[349]), .op(N742_t2) );
fim FAN_N742_3 ( .fault(fault), .net(N742), .FEN(FEN[350]), .op(N742_t3) );
fim FAN_N742_4 ( .fault(fault), .net(N742), .FEN(FEN[351]), .op(N742_t4) );
fim FAN_N599_0 ( .fault(fault), .net(N599), .FEN(FEN[352]), .op(N599_t0) );
fim FAN_N599_1 ( .fault(fault), .net(N599), .FEN(FEN[353]), .op(N599_t1) );
fim FAN_N599_2 ( .fault(fault), .net(N599), .FEN(FEN[354]), .op(N599_t2) );
fim FAN_N599_3 ( .fault(fault), .net(N599), .FEN(FEN[355]), .op(N599_t3) );
fim FAN_N727_0 ( .fault(fault), .net(N727), .FEN(FEN[356]), .op(N727_t0) );
fim FAN_N727_1 ( .fault(fault), .net(N727), .FEN(FEN[357]), .op(N727_t1) );
fim FAN_N727_2 ( .fault(fault), .net(N727), .FEN(FEN[358]), .op(N727_t2) );
fim FAN_N727_3 ( .fault(fault), .net(N727), .FEN(FEN[359]), .op(N727_t3) );
fim FAN_N727_4 ( .fault(fault), .net(N727), .FEN(FEN[360]), .op(N727_t4) );
fim FAN_N721_0 ( .fault(fault), .net(N721), .FEN(FEN[361]), .op(N721_t0) );
fim FAN_N721_1 ( .fault(fault), .net(N721), .FEN(FEN[362]), .op(N721_t1) );
fim FAN_N721_2 ( .fault(fault), .net(N721), .FEN(FEN[363]), .op(N721_t2) );
fim FAN_N721_3 ( .fault(fault), .net(N721), .FEN(FEN[364]), .op(N721_t3) );
fim FAN_N721_4 ( .fault(fault), .net(N721), .FEN(FEN[365]), .op(N721_t4) );
fim FAN_N715_0 ( .fault(fault), .net(N715), .FEN(FEN[366]), .op(N715_t0) );
fim FAN_N715_1 ( .fault(fault), .net(N715), .FEN(FEN[367]), .op(N715_t1) );
fim FAN_N715_2 ( .fault(fault), .net(N715), .FEN(FEN[368]), .op(N715_t2) );
fim FAN_N715_3 ( .fault(fault), .net(N715), .FEN(FEN[369]), .op(N715_t3) );
fim FAN_N715_4 ( .fault(fault), .net(N715), .FEN(FEN[370]), .op(N715_t4) );
fim FAN_N734_0 ( .fault(fault), .net(N734), .FEN(FEN[371]), .op(N734_t0) );
fim FAN_N734_1 ( .fault(fault), .net(N734), .FEN(FEN[372]), .op(N734_t1) );
fim FAN_N734_2 ( .fault(fault), .net(N734), .FEN(FEN[373]), .op(N734_t2) );
fim FAN_N734_3 ( .fault(fault), .net(N734), .FEN(FEN[374]), .op(N734_t3) );
fim FAN_N734_4 ( .fault(fault), .net(N734), .FEN(FEN[375]), .op(N734_t4) );
fim FAN_N734_5 ( .fault(fault), .net(N734), .FEN(FEN[376]), .op(N734_t5) );
fim FAN_N734_6 ( .fault(fault), .net(N734), .FEN(FEN[377]), .op(N734_t6) );
fim FAN_N708_0 ( .fault(fault), .net(N708), .FEN(FEN[378]), .op(N708_t0) );
fim FAN_N708_1 ( .fault(fault), .net(N708), .FEN(FEN[379]), .op(N708_t1) );
fim FAN_N708_2 ( .fault(fault), .net(N708), .FEN(FEN[380]), .op(N708_t2) );
fim FAN_N708_3 ( .fault(fault), .net(N708), .FEN(FEN[381]), .op(N708_t3) );
fim FAN_N708_4 ( .fault(fault), .net(N708), .FEN(FEN[382]), .op(N708_t4) );
fim FAN_N708_5 ( .fault(fault), .net(N708), .FEN(FEN[383]), .op(N708_t5) );
fim FAN_N806_0 ( .fault(fault), .net(N806), .FEN(FEN[384]), .op(N806_t0) );
fim FAN_N806_1 ( .fault(fault), .net(N806), .FEN(FEN[385]), .op(N806_t1) );
fim FAN_N806_2 ( .fault(fault), .net(N806), .FEN(FEN[386]), .op(N806_t2) );
fim FAN_N806_3 ( .fault(fault), .net(N806), .FEN(FEN[387]), .op(N806_t3) );
fim FAN_N806_4 ( .fault(fault), .net(N806), .FEN(FEN[388]), .op(N806_t4) );
fim FAN_N800_0 ( .fault(fault), .net(N800), .FEN(FEN[389]), .op(N800_t0) );
fim FAN_N800_1 ( .fault(fault), .net(N800), .FEN(FEN[390]), .op(N800_t1) );
fim FAN_N800_2 ( .fault(fault), .net(N800), .FEN(FEN[391]), .op(N800_t2) );
fim FAN_N800_3 ( .fault(fault), .net(N800), .FEN(FEN[392]), .op(N800_t3) );
fim FAN_N800_4 ( .fault(fault), .net(N800), .FEN(FEN[393]), .op(N800_t4) );
fim FAN_N794_0 ( .fault(fault), .net(N794), .FEN(FEN[394]), .op(N794_t0) );
fim FAN_N794_1 ( .fault(fault), .net(N794), .FEN(FEN[395]), .op(N794_t1) );
fim FAN_N794_2 ( .fault(fault), .net(N794), .FEN(FEN[396]), .op(N794_t2) );
fim FAN_N794_3 ( .fault(fault), .net(N794), .FEN(FEN[397]), .op(N794_t3) );
fim FAN_N794_4 ( .fault(fault), .net(N794), .FEN(FEN[398]), .op(N794_t4) );
fim FAN_N786_0 ( .fault(fault), .net(N786), .FEN(FEN[399]), .op(N786_t0) );
fim FAN_N786_1 ( .fault(fault), .net(N786), .FEN(FEN[400]), .op(N786_t1) );
fim FAN_N786_2 ( .fault(fault), .net(N786), .FEN(FEN[401]), .op(N786_t2) );
fim FAN_N786_3 ( .fault(fault), .net(N786), .FEN(FEN[402]), .op(N786_t3) );
fim FAN_N786_4 ( .fault(fault), .net(N786), .FEN(FEN[403]), .op(N786_t4) );
fim FAN_N786_5 ( .fault(fault), .net(N786), .FEN(FEN[404]), .op(N786_t5) );
fim FAN_N786_6 ( .fault(fault), .net(N786), .FEN(FEN[405]), .op(N786_t6) );
fim FAN_N780_0 ( .fault(fault), .net(N780), .FEN(FEN[406]), .op(N780_t0) );
fim FAN_N780_1 ( .fault(fault), .net(N780), .FEN(FEN[407]), .op(N780_t1) );
fim FAN_N780_2 ( .fault(fault), .net(N780), .FEN(FEN[408]), .op(N780_t2) );
fim FAN_N780_3 ( .fault(fault), .net(N780), .FEN(FEN[409]), .op(N780_t3) );
fim FAN_N780_4 ( .fault(fault), .net(N780), .FEN(FEN[410]), .op(N780_t4) );
fim FAN_N774_0 ( .fault(fault), .net(N774), .FEN(FEN[411]), .op(N774_t0) );
fim FAN_N774_1 ( .fault(fault), .net(N774), .FEN(FEN[412]), .op(N774_t1) );
fim FAN_N774_2 ( .fault(fault), .net(N774), .FEN(FEN[413]), .op(N774_t2) );
fim FAN_N774_3 ( .fault(fault), .net(N774), .FEN(FEN[414]), .op(N774_t3) );
fim FAN_N774_4 ( .fault(fault), .net(N774), .FEN(FEN[415]), .op(N774_t4) );
fim FAN_N768_0 ( .fault(fault), .net(N768), .FEN(FEN[416]), .op(N768_t0) );
fim FAN_N768_1 ( .fault(fault), .net(N768), .FEN(FEN[417]), .op(N768_t1) );
fim FAN_N768_2 ( .fault(fault), .net(N768), .FEN(FEN[418]), .op(N768_t2) );
fim FAN_N768_3 ( .fault(fault), .net(N768), .FEN(FEN[419]), .op(N768_t3) );
fim FAN_N768_4 ( .fault(fault), .net(N768), .FEN(FEN[420]), .op(N768_t4) );
fim FAN_N762_0 ( .fault(fault), .net(N762), .FEN(FEN[421]), .op(N762_t0) );
fim FAN_N762_1 ( .fault(fault), .net(N762), .FEN(FEN[422]), .op(N762_t1) );
fim FAN_N762_2 ( .fault(fault), .net(N762), .FEN(FEN[423]), .op(N762_t2) );
fim FAN_N762_3 ( .fault(fault), .net(N762), .FEN(FEN[424]), .op(N762_t3) );
fim FAN_N762_4 ( .fault(fault), .net(N762), .FEN(FEN[425]), .op(N762_t4) );
fim FAN_N636_0 ( .fault(fault), .net(N636), .FEN(FEN[426]), .op(N636_t0) );
fim FAN_N636_1 ( .fault(fault), .net(N636), .FEN(FEN[427]), .op(N636_t1) );
fim FAN_N636_2 ( .fault(fault), .net(N636), .FEN(FEN[428]), .op(N636_t2) );
fim FAN_N636_3 ( .fault(fault), .net(N636), .FEN(FEN[429]), .op(N636_t3) );
fim FAN_N865_0 ( .fault(fault), .net(N865), .FEN(FEN[430]), .op(N865_t0) );
fim FAN_N865_1 ( .fault(fault), .net(N865), .FEN(FEN[431]), .op(N865_t1) );
fim FAN_N865_2 ( .fault(fault), .net(N865), .FEN(FEN[432]), .op(N865_t2) );
fim FAN_N865_3 ( .fault(fault), .net(N865), .FEN(FEN[433]), .op(N865_t3) );
fim FAN_N865_4 ( .fault(fault), .net(N865), .FEN(FEN[434]), .op(N865_t4) );
fim FAN_N859_0 ( .fault(fault), .net(N859), .FEN(FEN[435]), .op(N859_t0) );
fim FAN_N859_1 ( .fault(fault), .net(N859), .FEN(FEN[436]), .op(N859_t1) );
fim FAN_N859_2 ( .fault(fault), .net(N859), .FEN(FEN[437]), .op(N859_t2) );
fim FAN_N859_3 ( .fault(fault), .net(N859), .FEN(FEN[438]), .op(N859_t3) );
fim FAN_N859_4 ( .fault(fault), .net(N859), .FEN(FEN[439]), .op(N859_t4) );
fim FAN_N853_0 ( .fault(fault), .net(N853), .FEN(FEN[440]), .op(N853_t0) );
fim FAN_N853_1 ( .fault(fault), .net(N853), .FEN(FEN[441]), .op(N853_t1) );
fim FAN_N853_2 ( .fault(fault), .net(N853), .FEN(FEN[442]), .op(N853_t2) );
fim FAN_N853_3 ( .fault(fault), .net(N853), .FEN(FEN[443]), .op(N853_t3) );
fim FAN_N853_4 ( .fault(fault), .net(N853), .FEN(FEN[444]), .op(N853_t4) );
fim FAN_N845_0 ( .fault(fault), .net(N845), .FEN(FEN[445]), .op(N845_t0) );
fim FAN_N845_1 ( .fault(fault), .net(N845), .FEN(FEN[446]), .op(N845_t1) );
fim FAN_N845_2 ( .fault(fault), .net(N845), .FEN(FEN[447]), .op(N845_t2) );
fim FAN_N845_3 ( .fault(fault), .net(N845), .FEN(FEN[448]), .op(N845_t3) );
fim FAN_N845_4 ( .fault(fault), .net(N845), .FEN(FEN[449]), .op(N845_t4) );
fim FAN_N845_5 ( .fault(fault), .net(N845), .FEN(FEN[450]), .op(N845_t5) );
fim FAN_N845_6 ( .fault(fault), .net(N845), .FEN(FEN[451]), .op(N845_t6) );
fim FAN_N839_0 ( .fault(fault), .net(N839), .FEN(FEN[452]), .op(N839_t0) );
fim FAN_N839_1 ( .fault(fault), .net(N839), .FEN(FEN[453]), .op(N839_t1) );
fim FAN_N839_2 ( .fault(fault), .net(N839), .FEN(FEN[454]), .op(N839_t2) );
fim FAN_N839_3 ( .fault(fault), .net(N839), .FEN(FEN[455]), .op(N839_t3) );
fim FAN_N839_4 ( .fault(fault), .net(N839), .FEN(FEN[456]), .op(N839_t4) );
fim FAN_N833_0 ( .fault(fault), .net(N833), .FEN(FEN[457]), .op(N833_t0) );
fim FAN_N833_1 ( .fault(fault), .net(N833), .FEN(FEN[458]), .op(N833_t1) );
fim FAN_N833_2 ( .fault(fault), .net(N833), .FEN(FEN[459]), .op(N833_t2) );
fim FAN_N833_3 ( .fault(fault), .net(N833), .FEN(FEN[460]), .op(N833_t3) );
fim FAN_N833_4 ( .fault(fault), .net(N833), .FEN(FEN[461]), .op(N833_t4) );
fim FAN_N827_0 ( .fault(fault), .net(N827), .FEN(FEN[462]), .op(N827_t0) );
fim FAN_N827_1 ( .fault(fault), .net(N827), .FEN(FEN[463]), .op(N827_t1) );
fim FAN_N827_2 ( .fault(fault), .net(N827), .FEN(FEN[464]), .op(N827_t2) );
fim FAN_N827_3 ( .fault(fault), .net(N827), .FEN(FEN[465]), .op(N827_t3) );
fim FAN_N827_4 ( .fault(fault), .net(N827), .FEN(FEN[466]), .op(N827_t4) );
fim FAN_N821_0 ( .fault(fault), .net(N821), .FEN(FEN[467]), .op(N821_t0) );
fim FAN_N821_1 ( .fault(fault), .net(N821), .FEN(FEN[468]), .op(N821_t1) );
fim FAN_N821_2 ( .fault(fault), .net(N821), .FEN(FEN[469]), .op(N821_t2) );
fim FAN_N821_3 ( .fault(fault), .net(N821), .FEN(FEN[470]), .op(N821_t3) );
fim FAN_N821_4 ( .fault(fault), .net(N821), .FEN(FEN[471]), .op(N821_t4) );
fim FAN_N814_0 ( .fault(fault), .net(N814), .FEN(FEN[472]), .op(N814_t0) );
fim FAN_N814_1 ( .fault(fault), .net(N814), .FEN(FEN[473]), .op(N814_t1) );
fim FAN_N814_2 ( .fault(fault), .net(N814), .FEN(FEN[474]), .op(N814_t2) );
fim FAN_N814_3 ( .fault(fault), .net(N814), .FEN(FEN[475]), .op(N814_t3) );
fim FAN_N814_4 ( .fault(fault), .net(N814), .FEN(FEN[476]), .op(N814_t4) );
fim FAN_N814_5 ( .fault(fault), .net(N814), .FEN(FEN[477]), .op(N814_t5) );
fim FAN_N1116_0 ( .fault(fault), .net(N1116), .FEN(FEN[478]), .op(N1116_t0) );
fim FAN_N1116_1 ( .fault(fault), .net(N1116), .FEN(FEN[479]), .op(N1116_t1) );
fim FAN_N957_0 ( .fault(fault), .net(N957), .FEN(FEN[480]), .op(N957_t0) );
fim FAN_N957_1 ( .fault(fault), .net(N957), .FEN(FEN[481]), .op(N957_t1) );
fim FAN_N957_2 ( .fault(fault), .net(N957), .FEN(FEN[482]), .op(N957_t2) );
fim FAN_N957_3 ( .fault(fault), .net(N957), .FEN(FEN[483]), .op(N957_t3) );
fim FAN_N957_4 ( .fault(fault), .net(N957), .FEN(FEN[484]), .op(N957_t4) );
fim FAN_N957_5 ( .fault(fault), .net(N957), .FEN(FEN[485]), .op(N957_t5) );
fim FAN_N1029_0 ( .fault(fault), .net(N1029), .FEN(FEN[486]), .op(N1029_t0) );
fim FAN_N1029_1 ( .fault(fault), .net(N1029), .FEN(FEN[487]), .op(N1029_t1) );
fim FAN_N1125_0 ( .fault(fault), .net(N1125), .FEN(FEN[488]), .op(N1125_t0) );
fim FAN_N1125_1 ( .fault(fault), .net(N1125), .FEN(FEN[489]), .op(N1125_t1) );
fim FAN_N1125_2 ( .fault(fault), .net(N1125), .FEN(FEN[490]), .op(N1125_t2) );
fim FAN_N1125_3 ( .fault(fault), .net(N1125), .FEN(FEN[491]), .op(N1125_t3) );
fim FAN_N1125_4 ( .fault(fault), .net(N1125), .FEN(FEN[492]), .op(N1125_t4) );
fim FAN_N1125_5 ( .fault(fault), .net(N1125), .FEN(FEN[493]), .op(N1125_t5) );
fim FAN_N1136_0 ( .fault(fault), .net(N1136), .FEN(FEN[494]), .op(N1136_t0) );
fim FAN_N1136_1 ( .fault(fault), .net(N1136), .FEN(FEN[495]), .op(N1136_t1) );
fim FAN_N1136_2 ( .fault(fault), .net(N1136), .FEN(FEN[496]), .op(N1136_t2) );
fim FAN_N1136_3 ( .fault(fault), .net(N1136), .FEN(FEN[497]), .op(N1136_t3) );
fim FAN_N1147_0 ( .fault(fault), .net(N1147), .FEN(FEN[498]), .op(N1147_t0) );
fim FAN_N1147_1 ( .fault(fault), .net(N1147), .FEN(FEN[499]), .op(N1147_t1) );
fim FAN_N1147_2 ( .fault(fault), .net(N1147), .FEN(FEN[500]), .op(N1147_t2) );
fim FAN_N1147_3 ( .fault(fault), .net(N1147), .FEN(FEN[501]), .op(N1147_t3) );
fim FAN_N1147_4 ( .fault(fault), .net(N1147), .FEN(FEN[502]), .op(N1147_t4) );
fim FAN_N1147_5 ( .fault(fault), .net(N1147), .FEN(FEN[503]), .op(N1147_t5) );
fim FAN_N1160_0 ( .fault(fault), .net(N1160), .FEN(FEN[504]), .op(N1160_t0) );
fim FAN_N1160_1 ( .fault(fault), .net(N1160), .FEN(FEN[505]), .op(N1160_t1) );
fim FAN_N1160_2 ( .fault(fault), .net(N1160), .FEN(FEN[506]), .op(N1160_t2) );
fim FAN_N1160_3 ( .fault(fault), .net(N1160), .FEN(FEN[507]), .op(N1160_t3) );
fim FAN_N1160_4 ( .fault(fault), .net(N1160), .FEN(FEN[508]), .op(N1160_t4) );
fim FAN_N1160_5 ( .fault(fault), .net(N1160), .FEN(FEN[509]), .op(N1160_t5) );
fim FAN_N1284_0 ( .fault(fault), .net(N1284), .FEN(FEN[510]), .op(N1284_t0) );
fim FAN_N1284_1 ( .fault(fault), .net(N1284), .FEN(FEN[511]), .op(N1284_t1) );
fim FAN_N1287_0 ( .fault(fault), .net(N1287), .FEN(FEN[512]), .op(N1287_t0) );
fim FAN_N1287_1 ( .fault(fault), .net(N1287), .FEN(FEN[513]), .op(N1287_t1) );
fim FAN_N1290_0 ( .fault(fault), .net(N1290), .FEN(FEN[514]), .op(N1290_t0) );
fim FAN_N1290_1 ( .fault(fault), .net(N1290), .FEN(FEN[515]), .op(N1290_t1) );
fim FAN_N1293_0 ( .fault(fault), .net(N1293), .FEN(FEN[516]), .op(N1293_t0) );
fim FAN_N1293_1 ( .fault(fault), .net(N1293), .FEN(FEN[517]), .op(N1293_t1) );
fim FAN_N1296_0 ( .fault(fault), .net(N1296), .FEN(FEN[518]), .op(N1296_t0) );
fim FAN_N1296_1 ( .fault(fault), .net(N1296), .FEN(FEN[519]), .op(N1296_t1) );
fim FAN_N1299_0 ( .fault(fault), .net(N1299), .FEN(FEN[520]), .op(N1299_t0) );
fim FAN_N1299_1 ( .fault(fault), .net(N1299), .FEN(FEN[521]), .op(N1299_t1) );
fim FAN_N1302_0 ( .fault(fault), .net(N1302), .FEN(FEN[522]), .op(N1302_t0) );
fim FAN_N1302_1 ( .fault(fault), .net(N1302), .FEN(FEN[523]), .op(N1302_t1) );
fim FAN_N1305_0 ( .fault(fault), .net(N1305), .FEN(FEN[524]), .op(N1305_t0) );
fim FAN_N1305_1 ( .fault(fault), .net(N1305), .FEN(FEN[525]), .op(N1305_t1) );
fim FAN_N1308_0 ( .fault(fault), .net(N1308), .FEN(FEN[526]), .op(N1308_t0) );
fim FAN_N1308_1 ( .fault(fault), .net(N1308), .FEN(FEN[527]), .op(N1308_t1) );
fim FAN_N1311_0 ( .fault(fault), .net(N1311), .FEN(FEN[528]), .op(N1311_t0) );
fim FAN_N1311_1 ( .fault(fault), .net(N1311), .FEN(FEN[529]), .op(N1311_t1) );
fim FAN_N1314_0 ( .fault(fault), .net(N1314), .FEN(FEN[530]), .op(N1314_t0) );
fim FAN_N1314_1 ( .fault(fault), .net(N1314), .FEN(FEN[531]), .op(N1314_t1) );
fim FAN_N1317_0 ( .fault(fault), .net(N1317), .FEN(FEN[532]), .op(N1317_t0) );
fim FAN_N1317_1 ( .fault(fault), .net(N1317), .FEN(FEN[533]), .op(N1317_t1) );
fim FAN_N1320_0 ( .fault(fault), .net(N1320), .FEN(FEN[534]), .op(N1320_t0) );
fim FAN_N1320_1 ( .fault(fault), .net(N1320), .FEN(FEN[535]), .op(N1320_t1) );
fim FAN_N1323_0 ( .fault(fault), .net(N1323), .FEN(FEN[536]), .op(N1323_t0) );
fim FAN_N1323_1 ( .fault(fault), .net(N1323), .FEN(FEN[537]), .op(N1323_t1) );
fim FAN_N1175_0 ( .fault(fault), .net(N1175), .FEN(FEN[538]), .op(N1175_t0) );
fim FAN_N1175_1 ( .fault(fault), .net(N1175), .FEN(FEN[539]), .op(N1175_t1) );
fim FAN_N1175_2 ( .fault(fault), .net(N1175), .FEN(FEN[540]), .op(N1175_t2) );
fim FAN_N1175_3 ( .fault(fault), .net(N1175), .FEN(FEN[541]), .op(N1175_t3) );
fim FAN_N1175_4 ( .fault(fault), .net(N1175), .FEN(FEN[542]), .op(N1175_t4) );
fim FAN_N1175_5 ( .fault(fault), .net(N1175), .FEN(FEN[543]), .op(N1175_t5) );
fim FAN_N1182_0 ( .fault(fault), .net(N1182), .FEN(FEN[544]), .op(N1182_t0) );
fim FAN_N1182_1 ( .fault(fault), .net(N1182), .FEN(FEN[545]), .op(N1182_t1) );
fim FAN_N1182_2 ( .fault(fault), .net(N1182), .FEN(FEN[546]), .op(N1182_t2) );
fim FAN_N1182_3 ( .fault(fault), .net(N1182), .FEN(FEN[547]), .op(N1182_t3) );
fim FAN_N1182_4 ( .fault(fault), .net(N1182), .FEN(FEN[548]), .op(N1182_t4) );
fim FAN_N1182_5 ( .fault(fault), .net(N1182), .FEN(FEN[549]), .op(N1182_t5) );
fim FAN_N1326_0 ( .fault(fault), .net(N1326), .FEN(FEN[550]), .op(N1326_t0) );
fim FAN_N1326_1 ( .fault(fault), .net(N1326), .FEN(FEN[551]), .op(N1326_t1) );
fim FAN_N1329_0 ( .fault(fault), .net(N1329), .FEN(FEN[552]), .op(N1329_t0) );
fim FAN_N1329_1 ( .fault(fault), .net(N1329), .FEN(FEN[553]), .op(N1329_t1) );
fim FAN_N1332_0 ( .fault(fault), .net(N1332), .FEN(FEN[554]), .op(N1332_t0) );
fim FAN_N1332_1 ( .fault(fault), .net(N1332), .FEN(FEN[555]), .op(N1332_t1) );
fim FAN_N1335_0 ( .fault(fault), .net(N1335), .FEN(FEN[556]), .op(N1335_t0) );
fim FAN_N1335_1 ( .fault(fault), .net(N1335), .FEN(FEN[557]), .op(N1335_t1) );
fim FAN_N1338_0 ( .fault(fault), .net(N1338), .FEN(FEN[558]), .op(N1338_t0) );
fim FAN_N1338_1 ( .fault(fault), .net(N1338), .FEN(FEN[559]), .op(N1338_t1) );
fim FAN_N1341_0 ( .fault(fault), .net(N1341), .FEN(FEN[560]), .op(N1341_t0) );
fim FAN_N1341_1 ( .fault(fault), .net(N1341), .FEN(FEN[561]), .op(N1341_t1) );
fim FAN_N1344_0 ( .fault(fault), .net(N1344), .FEN(FEN[562]), .op(N1344_t0) );
fim FAN_N1344_1 ( .fault(fault), .net(N1344), .FEN(FEN[563]), .op(N1344_t1) );
fim FAN_N1347_0 ( .fault(fault), .net(N1347), .FEN(FEN[564]), .op(N1347_t0) );
fim FAN_N1347_1 ( .fault(fault), .net(N1347), .FEN(FEN[565]), .op(N1347_t1) );
fim FAN_N1350_0 ( .fault(fault), .net(N1350), .FEN(FEN[566]), .op(N1350_t0) );
fim FAN_N1350_1 ( .fault(fault), .net(N1350), .FEN(FEN[567]), .op(N1350_t1) );
fim FAN_N1353_0 ( .fault(fault), .net(N1353), .FEN(FEN[568]), .op(N1353_t0) );
fim FAN_N1353_1 ( .fault(fault), .net(N1353), .FEN(FEN[569]), .op(N1353_t1) );
fim FAN_N1356_0 ( .fault(fault), .net(N1356), .FEN(FEN[570]), .op(N1356_t0) );
fim FAN_N1356_1 ( .fault(fault), .net(N1356), .FEN(FEN[571]), .op(N1356_t1) );
fim FAN_N1359_0 ( .fault(fault), .net(N1359), .FEN(FEN[572]), .op(N1359_t0) );
fim FAN_N1359_1 ( .fault(fault), .net(N1359), .FEN(FEN[573]), .op(N1359_t1) );
fim FAN_N1362_0 ( .fault(fault), .net(N1362), .FEN(FEN[574]), .op(N1362_t0) );
fim FAN_N1362_1 ( .fault(fault), .net(N1362), .FEN(FEN[575]), .op(N1362_t1) );
fim FAN_N1365_0 ( .fault(fault), .net(N1365), .FEN(FEN[576]), .op(N1365_t0) );
fim FAN_N1365_1 ( .fault(fault), .net(N1365), .FEN(FEN[577]), .op(N1365_t1) );
fim FAN_N1368_0 ( .fault(fault), .net(N1368), .FEN(FEN[578]), .op(N1368_t0) );
fim FAN_N1368_1 ( .fault(fault), .net(N1368), .FEN(FEN[579]), .op(N1368_t1) );
fim FAN_N1371_0 ( .fault(fault), .net(N1371), .FEN(FEN[580]), .op(N1371_t0) );
fim FAN_N1371_1 ( .fault(fault), .net(N1371), .FEN(FEN[581]), .op(N1371_t1) );
fim FAN_N1374_0 ( .fault(fault), .net(N1374), .FEN(FEN[582]), .op(N1374_t0) );
fim FAN_N1374_1 ( .fault(fault), .net(N1374), .FEN(FEN[583]), .op(N1374_t1) );
fim FAN_N1377_0 ( .fault(fault), .net(N1377), .FEN(FEN[584]), .op(N1377_t0) );
fim FAN_N1377_1 ( .fault(fault), .net(N1377), .FEN(FEN[585]), .op(N1377_t1) );
fim FAN_N1199_0 ( .fault(fault), .net(N1199), .FEN(FEN[586]), .op(N1199_t0) );
fim FAN_N1199_1 ( .fault(fault), .net(N1199), .FEN(FEN[587]), .op(N1199_t1) );
fim FAN_N1194_0 ( .fault(fault), .net(N1194), .FEN(FEN[588]), .op(N1194_t0) );
fim FAN_N1194_1 ( .fault(fault), .net(N1194), .FEN(FEN[589]), .op(N1194_t1) );
fim FAN_N1194_2 ( .fault(fault), .net(N1194), .FEN(FEN[590]), .op(N1194_t2) );
fim FAN_N1194_3 ( .fault(fault), .net(N1194), .FEN(FEN[591]), .op(N1194_t3) );
fim FAN_N1211_0 ( .fault(fault), .net(N1211), .FEN(FEN[592]), .op(N1211_t0) );
fim FAN_N1211_1 ( .fault(fault), .net(N1211), .FEN(FEN[593]), .op(N1211_t1) );
fim FAN_N1211_2 ( .fault(fault), .net(N1211), .FEN(FEN[594]), .op(N1211_t2) );
fim FAN_N1211_3 ( .fault(fault), .net(N1211), .FEN(FEN[595]), .op(N1211_t3) );
fim FAN_N1211_4 ( .fault(fault), .net(N1211), .FEN(FEN[596]), .op(N1211_t4) );
fim FAN_N1211_5 ( .fault(fault), .net(N1211), .FEN(FEN[597]), .op(N1211_t5) );
fim FAN_N44_0 ( .fault(fault), .net(N44), .FEN(FEN[598]), .op(N44_t0) );
fim FAN_N44_1 ( .fault(fault), .net(N44), .FEN(FEN[599]), .op(N44_t1) );
fim FAN_N41_0 ( .fault(fault), .net(N41), .FEN(FEN[600]), .op(N41_t0) );
fim FAN_N41_1 ( .fault(fault), .net(N41), .FEN(FEN[601]), .op(N41_t1) );
fim FAN_N29_0 ( .fault(fault), .net(N29), .FEN(FEN[602]), .op(N29_t0) );
fim FAN_N29_1 ( .fault(fault), .net(N29), .FEN(FEN[603]), .op(N29_t1) );
fim FAN_N26_0 ( .fault(fault), .net(N26), .FEN(FEN[604]), .op(N26_t0) );
fim FAN_N26_1 ( .fault(fault), .net(N26), .FEN(FEN[605]), .op(N26_t1) );
fim FAN_N23_0 ( .fault(fault), .net(N23), .FEN(FEN[606]), .op(N23_t0) );
fim FAN_N23_1 ( .fault(fault), .net(N23), .FEN(FEN[607]), .op(N23_t1) );
fim FAN_N1380_0 ( .fault(fault), .net(N1380), .FEN(FEN[608]), .op(N1380_t0) );
fim FAN_N1380_1 ( .fault(fault), .net(N1380), .FEN(FEN[609]), .op(N1380_t1) );
fim FAN_N1383_0 ( .fault(fault), .net(N1383), .FEN(FEN[610]), .op(N1383_t0) );
fim FAN_N1383_1 ( .fault(fault), .net(N1383), .FEN(FEN[611]), .op(N1383_t1) );
fim FAN_N1386_0 ( .fault(fault), .net(N1386), .FEN(FEN[612]), .op(N1386_t0) );
fim FAN_N1386_1 ( .fault(fault), .net(N1386), .FEN(FEN[613]), .op(N1386_t1) );
fim FAN_N1389_0 ( .fault(fault), .net(N1389), .FEN(FEN[614]), .op(N1389_t0) );
fim FAN_N1389_1 ( .fault(fault), .net(N1389), .FEN(FEN[615]), .op(N1389_t1) );
fim FAN_N1392_0 ( .fault(fault), .net(N1392), .FEN(FEN[616]), .op(N1392_t0) );
fim FAN_N1392_1 ( .fault(fault), .net(N1392), .FEN(FEN[617]), .op(N1392_t1) );
fim FAN_N1395_0 ( .fault(fault), .net(N1395), .FEN(FEN[618]), .op(N1395_t0) );
fim FAN_N1395_1 ( .fault(fault), .net(N1395), .FEN(FEN[619]), .op(N1395_t1) );
fim FAN_N1398_0 ( .fault(fault), .net(N1398), .FEN(FEN[620]), .op(N1398_t0) );
fim FAN_N1398_1 ( .fault(fault), .net(N1398), .FEN(FEN[621]), .op(N1398_t1) );
fim FAN_N1401_0 ( .fault(fault), .net(N1401), .FEN(FEN[622]), .op(N1401_t0) );
fim FAN_N1401_1 ( .fault(fault), .net(N1401), .FEN(FEN[623]), .op(N1401_t1) );
fim FAN_N1404_0 ( .fault(fault), .net(N1404), .FEN(FEN[624]), .op(N1404_t0) );
fim FAN_N1404_1 ( .fault(fault), .net(N1404), .FEN(FEN[625]), .op(N1404_t1) );
fim FAN_N1407_0 ( .fault(fault), .net(N1407), .FEN(FEN[626]), .op(N1407_t0) );
fim FAN_N1407_1 ( .fault(fault), .net(N1407), .FEN(FEN[627]), .op(N1407_t1) );
fim FAN_N1410_0 ( .fault(fault), .net(N1410), .FEN(FEN[628]), .op(N1410_t0) );
fim FAN_N1410_1 ( .fault(fault), .net(N1410), .FEN(FEN[629]), .op(N1410_t1) );
fim FAN_N1413_0 ( .fault(fault), .net(N1413), .FEN(FEN[630]), .op(N1413_t0) );
fim FAN_N1413_1 ( .fault(fault), .net(N1413), .FEN(FEN[631]), .op(N1413_t1) );
fim FAN_N1416_0 ( .fault(fault), .net(N1416), .FEN(FEN[632]), .op(N1416_t0) );
fim FAN_N1416_1 ( .fault(fault), .net(N1416), .FEN(FEN[633]), .op(N1416_t1) );
fim FAN_N1419_0 ( .fault(fault), .net(N1419), .FEN(FEN[634]), .op(N1419_t0) );
fim FAN_N1419_1 ( .fault(fault), .net(N1419), .FEN(FEN[635]), .op(N1419_t1) );
fim FAN_N1422_0 ( .fault(fault), .net(N1422), .FEN(FEN[636]), .op(N1422_t0) );
fim FAN_N1422_1 ( .fault(fault), .net(N1422), .FEN(FEN[637]), .op(N1422_t1) );
fim FAN_N1425_0 ( .fault(fault), .net(N1425), .FEN(FEN[638]), .op(N1425_t0) );
fim FAN_N1425_1 ( .fault(fault), .net(N1425), .FEN(FEN[639]), .op(N1425_t1) );
fim FAN_N1233_0 ( .fault(fault), .net(N1233), .FEN(FEN[640]), .op(N1233_t0) );
fim FAN_N1233_1 ( .fault(fault), .net(N1233), .FEN(FEN[641]), .op(N1233_t1) );
fim FAN_N1233_2 ( .fault(fault), .net(N1233), .FEN(FEN[642]), .op(N1233_t2) );
fim FAN_N1233_3 ( .fault(fault), .net(N1233), .FEN(FEN[643]), .op(N1233_t3) );
fim FAN_N1233_4 ( .fault(fault), .net(N1233), .FEN(FEN[644]), .op(N1233_t4) );
fim FAN_N1233_5 ( .fault(fault), .net(N1233), .FEN(FEN[645]), .op(N1233_t5) );
fim FAN_N1244_0 ( .fault(fault), .net(N1244), .FEN(FEN[646]), .op(N1244_t0) );
fim FAN_N1244_1 ( .fault(fault), .net(N1244), .FEN(FEN[647]), .op(N1244_t1) );
fim FAN_N1244_2 ( .fault(fault), .net(N1244), .FEN(FEN[648]), .op(N1244_t2) );
fim FAN_N1244_3 ( .fault(fault), .net(N1244), .FEN(FEN[649]), .op(N1244_t3) );
fim FAN_N1428_0 ( .fault(fault), .net(N1428), .FEN(FEN[650]), .op(N1428_t0) );
fim FAN_N1428_1 ( .fault(fault), .net(N1428), .FEN(FEN[651]), .op(N1428_t1) );
fim FAN_N1222_0 ( .fault(fault), .net(N1222), .FEN(FEN[652]), .op(N1222_t0) );
fim FAN_N1222_1 ( .fault(fault), .net(N1222), .FEN(FEN[653]), .op(N1222_t1) );
fim FAN_N1431_0 ( .fault(fault), .net(N1431), .FEN(FEN[654]), .op(N1431_t0) );
fim FAN_N1431_1 ( .fault(fault), .net(N1431), .FEN(FEN[655]), .op(N1431_t1) );
fim FAN_N1434_0 ( .fault(fault), .net(N1434), .FEN(FEN[656]), .op(N1434_t0) );
fim FAN_N1434_1 ( .fault(fault), .net(N1434), .FEN(FEN[657]), .op(N1434_t1) );
fim FAN_N1437_0 ( .fault(fault), .net(N1437), .FEN(FEN[658]), .op(N1437_t0) );
fim FAN_N1437_1 ( .fault(fault), .net(N1437), .FEN(FEN[659]), .op(N1437_t1) );
fim FAN_N1440_0 ( .fault(fault), .net(N1440), .FEN(FEN[660]), .op(N1440_t0) );
fim FAN_N1440_1 ( .fault(fault), .net(N1440), .FEN(FEN[661]), .op(N1440_t1) );
fim FAN_N1443_0 ( .fault(fault), .net(N1443), .FEN(FEN[662]), .op(N1443_t0) );
fim FAN_N1443_1 ( .fault(fault), .net(N1443), .FEN(FEN[663]), .op(N1443_t1) );
fim FAN_N1446_0 ( .fault(fault), .net(N1446), .FEN(FEN[664]), .op(N1446_t0) );
fim FAN_N1446_1 ( .fault(fault), .net(N1446), .FEN(FEN[665]), .op(N1446_t1) );
fim FAN_N1449_0 ( .fault(fault), .net(N1449), .FEN(FEN[666]), .op(N1449_t0) );
fim FAN_N1449_1 ( .fault(fault), .net(N1449), .FEN(FEN[667]), .op(N1449_t1) );
fim FAN_N1452_0 ( .fault(fault), .net(N1452), .FEN(FEN[668]), .op(N1452_t0) );
fim FAN_N1452_1 ( .fault(fault), .net(N1452), .FEN(FEN[669]), .op(N1452_t1) );
fim FAN_N1455_0 ( .fault(fault), .net(N1455), .FEN(FEN[670]), .op(N1455_t0) );
fim FAN_N1455_1 ( .fault(fault), .net(N1455), .FEN(FEN[671]), .op(N1455_t1) );
fim FAN_N1458_0 ( .fault(fault), .net(N1458), .FEN(FEN[672]), .op(N1458_t0) );
fim FAN_N1458_1 ( .fault(fault), .net(N1458), .FEN(FEN[673]), .op(N1458_t1) );
fim FAN_N1249_0 ( .fault(fault), .net(N1249), .FEN(FEN[674]), .op(N1249_t0) );
fim FAN_N1249_1 ( .fault(fault), .net(N1249), .FEN(FEN[675]), .op(N1249_t1) );
fim FAN_N1249_2 ( .fault(fault), .net(N1249), .FEN(FEN[676]), .op(N1249_t2) );
fim FAN_N1249_3 ( .fault(fault), .net(N1249), .FEN(FEN[677]), .op(N1249_t3) );
fim FAN_N1249_4 ( .fault(fault), .net(N1249), .FEN(FEN[678]), .op(N1249_t4) );
fim FAN_N1249_5 ( .fault(fault), .net(N1249), .FEN(FEN[679]), .op(N1249_t5) );
fim FAN_N1256_0 ( .fault(fault), .net(N1256), .FEN(FEN[680]), .op(N1256_t0) );
fim FAN_N1256_1 ( .fault(fault), .net(N1256), .FEN(FEN[681]), .op(N1256_t1) );
fim FAN_N1256_2 ( .fault(fault), .net(N1256), .FEN(FEN[682]), .op(N1256_t2) );
fim FAN_N1256_3 ( .fault(fault), .net(N1256), .FEN(FEN[683]), .op(N1256_t3) );
fim FAN_N1256_4 ( .fault(fault), .net(N1256), .FEN(FEN[684]), .op(N1256_t4) );
fim FAN_N1256_5 ( .fault(fault), .net(N1256), .FEN(FEN[685]), .op(N1256_t5) );
fim FAN_N1263_0 ( .fault(fault), .net(N1263), .FEN(FEN[686]), .op(N1263_t0) );
fim FAN_N1263_1 ( .fault(fault), .net(N1263), .FEN(FEN[687]), .op(N1263_t1) );
fim FAN_N1263_2 ( .fault(fault), .net(N1263), .FEN(FEN[688]), .op(N1263_t2) );
fim FAN_N1263_3 ( .fault(fault), .net(N1263), .FEN(FEN[689]), .op(N1263_t3) );
fim FAN_N1263_4 ( .fault(fault), .net(N1263), .FEN(FEN[690]), .op(N1263_t4) );
fim FAN_N1263_5 ( .fault(fault), .net(N1263), .FEN(FEN[691]), .op(N1263_t5) );
fim FAN_N47_0 ( .fault(fault), .net(N47), .FEN(FEN[692]), .op(N47_t0) );
fim FAN_N47_1 ( .fault(fault), .net(N47), .FEN(FEN[693]), .op(N47_t1) );
fim FAN_N35_0 ( .fault(fault), .net(N35), .FEN(FEN[694]), .op(N35_t0) );
fim FAN_N35_1 ( .fault(fault), .net(N35), .FEN(FEN[695]), .op(N35_t1) );
fim FAN_N32_0 ( .fault(fault), .net(N32), .FEN(FEN[696]), .op(N32_t0) );
fim FAN_N32_1 ( .fault(fault), .net(N32), .FEN(FEN[697]), .op(N32_t1) );
fim FAN_N50_0 ( .fault(fault), .net(N50), .FEN(FEN[698]), .op(N50_t0) );
fim FAN_N50_1 ( .fault(fault), .net(N50), .FEN(FEN[699]), .op(N50_t1) );
fim FAN_N66_0 ( .fault(fault), .net(N66), .FEN(FEN[700]), .op(N66_t0) );
fim FAN_N66_1 ( .fault(fault), .net(N66), .FEN(FEN[701]), .op(N66_t1) );
fim FAN_N1461_0 ( .fault(fault), .net(N1461), .FEN(FEN[702]), .op(N1461_t0) );
fim FAN_N1461_1 ( .fault(fault), .net(N1461), .FEN(FEN[703]), .op(N1461_t1) );
fim FAN_N1464_0 ( .fault(fault), .net(N1464), .FEN(FEN[704]), .op(N1464_t0) );
fim FAN_N1464_1 ( .fault(fault), .net(N1464), .FEN(FEN[705]), .op(N1464_t1) );
fim FAN_N1467_0 ( .fault(fault), .net(N1467), .FEN(FEN[706]), .op(N1467_t0) );
fim FAN_N1467_1 ( .fault(fault), .net(N1467), .FEN(FEN[707]), .op(N1467_t1) );
fim FAN_N1470_0 ( .fault(fault), .net(N1470), .FEN(FEN[708]), .op(N1470_t0) );
fim FAN_N1470_1 ( .fault(fault), .net(N1470), .FEN(FEN[709]), .op(N1470_t1) );
fim FAN_N1473_0 ( .fault(fault), .net(N1473), .FEN(FEN[710]), .op(N1473_t0) );
fim FAN_N1473_1 ( .fault(fault), .net(N1473), .FEN(FEN[711]), .op(N1473_t1) );
fim FAN_N1476_0 ( .fault(fault), .net(N1476), .FEN(FEN[712]), .op(N1476_t0) );
fim FAN_N1476_1 ( .fault(fault), .net(N1476), .FEN(FEN[713]), .op(N1476_t1) );
fim FAN_N1479_0 ( .fault(fault), .net(N1479), .FEN(FEN[714]), .op(N1479_t0) );
fim FAN_N1479_1 ( .fault(fault), .net(N1479), .FEN(FEN[715]), .op(N1479_t1) );
fim FAN_N1482_0 ( .fault(fault), .net(N1482), .FEN(FEN[716]), .op(N1482_t0) );
fim FAN_N1482_1 ( .fault(fault), .net(N1482), .FEN(FEN[717]), .op(N1482_t1) );
fim FAN_N1485_0 ( .fault(fault), .net(N1485), .FEN(FEN[718]), .op(N1485_t0) );
fim FAN_N1485_1 ( .fault(fault), .net(N1485), .FEN(FEN[719]), .op(N1485_t1) );
fim FAN_N1206_0 ( .fault(fault), .net(N1206), .FEN(FEN[720]), .op(N1206_t0) );
fim FAN_N1206_1 ( .fault(fault), .net(N1206), .FEN(FEN[721]), .op(N1206_t1) );
fim FAN_N1206_2 ( .fault(fault), .net(N1206), .FEN(FEN[722]), .op(N1206_t2) );
fim FAN_N1206_3 ( .fault(fault), .net(N1206), .FEN(FEN[723]), .op(N1206_t3) );
fim FAN_N1270_0 ( .fault(fault), .net(N1270), .FEN(FEN[724]), .op(N1270_t0) );
fim FAN_N1270_1 ( .fault(fault), .net(N1270), .FEN(FEN[725]), .op(N1270_t1) );
fim FAN_N1270_2 ( .fault(fault), .net(N1270), .FEN(FEN[726]), .op(N1270_t2) );
fim FAN_N1270_3 ( .fault(fault), .net(N1270), .FEN(FEN[727]), .op(N1270_t3) );
fim FAN_N1270_4 ( .fault(fault), .net(N1270), .FEN(FEN[728]), .op(N1270_t4) );
fim FAN_N1270_5 ( .fault(fault), .net(N1270), .FEN(FEN[729]), .op(N1270_t5) );
fim FAN_N1277_0 ( .fault(fault), .net(N1277), .FEN(FEN[730]), .op(N1277_t0) );
fim FAN_N1277_1 ( .fault(fault), .net(N1277), .FEN(FEN[731]), .op(N1277_t1) );
fim FAN_N1277_2 ( .fault(fault), .net(N1277), .FEN(FEN[732]), .op(N1277_t2) );
fim FAN_N1277_3 ( .fault(fault), .net(N1277), .FEN(FEN[733]), .op(N1277_t3) );
fim FAN_N1277_4 ( .fault(fault), .net(N1277), .FEN(FEN[734]), .op(N1277_t4) );
fim FAN_N1277_5 ( .fault(fault), .net(N1277), .FEN(FEN[735]), .op(N1277_t5) );
fim FAN_N1189_0 ( .fault(fault), .net(N1189), .FEN(FEN[736]), .op(N1189_t0) );
fim FAN_N1189_1 ( .fault(fault), .net(N1189), .FEN(FEN[737]), .op(N1189_t1) );
fim FAN_N1189_2 ( .fault(fault), .net(N1189), .FEN(FEN[738]), .op(N1189_t2) );
fim FAN_N1189_3 ( .fault(fault), .net(N1189), .FEN(FEN[739]), .op(N1189_t3) );
fim FAN_N1703_0 ( .fault(fault), .net(N1703), .FEN(FEN[740]), .op(N1703_t0) );
fim FAN_N1703_1 ( .fault(fault), .net(N1703), .FEN(FEN[741]), .op(N1703_t1) );
fim FAN_N1713_0 ( .fault(fault), .net(N1713), .FEN(FEN[742]), .op(N1713_t0) );
fim FAN_N1713_1 ( .fault(fault), .net(N1713), .FEN(FEN[743]), .op(N1713_t1) );
fim FAN_N1721_0 ( .fault(fault), .net(N1721), .FEN(FEN[744]), .op(N1721_t0) );
fim FAN_N1721_1 ( .fault(fault), .net(N1721), .FEN(FEN[745]), .op(N1721_t1) );
fim FAN_N1758_0 ( .fault(fault), .net(N1758), .FEN(FEN[746]), .op(N1758_t0) );
fim FAN_N1758_1 ( .fault(fault), .net(N1758), .FEN(FEN[747]), .op(N1758_t1) );
fim FAN_N1708_0 ( .fault(fault), .net(N1708), .FEN(FEN[748]), .op(N1708_t0) );
fim FAN_N1708_1 ( .fault(fault), .net(N1708), .FEN(FEN[749]), .op(N1708_t1) );
fim FAN_N1537_0 ( .fault(fault), .net(N1537), .FEN(FEN[750]), .op(N1537_t0) );
fim FAN_N1537_1 ( .fault(fault), .net(N1537), .FEN(FEN[751]), .op(N1537_t1) );
fim FAN_N1537_2 ( .fault(fault), .net(N1537), .FEN(FEN[752]), .op(N1537_t2) );
fim FAN_N1537_3 ( .fault(fault), .net(N1537), .FEN(FEN[753]), .op(N1537_t3) );
fim FAN_N1537_4 ( .fault(fault), .net(N1537), .FEN(FEN[754]), .op(N1537_t4) );
fim FAN_N1551_0 ( .fault(fault), .net(N1551), .FEN(FEN[755]), .op(N1551_t0) );
fim FAN_N1551_1 ( .fault(fault), .net(N1551), .FEN(FEN[756]), .op(N1551_t1) );
fim FAN_N1783_0 ( .fault(fault), .net(N1783), .FEN(FEN[757]), .op(N1783_t0) );
fim FAN_N1783_1 ( .fault(fault), .net(N1783), .FEN(FEN[758]), .op(N1783_t1) );
fim FAN_N1783_2 ( .fault(fault), .net(N1783), .FEN(FEN[759]), .op(N1783_t2) );
fim FAN_N1783_3 ( .fault(fault), .net(N1783), .FEN(FEN[760]), .op(N1783_t3) );
fim FAN_N1783_4 ( .fault(fault), .net(N1783), .FEN(FEN[761]), .op(N1783_t4) );
fim FAN_N1789_0 ( .fault(fault), .net(N1789), .FEN(FEN[762]), .op(N1789_t0) );
fim FAN_N1789_1 ( .fault(fault), .net(N1789), .FEN(FEN[763]), .op(N1789_t1) );
fim FAN_N1789_2 ( .fault(fault), .net(N1789), .FEN(FEN[764]), .op(N1789_t2) );
fim FAN_N1799_0 ( .fault(fault), .net(N1799), .FEN(FEN[765]), .op(N1799_t0) );
fim FAN_N1799_1 ( .fault(fault), .net(N1799), .FEN(FEN[766]), .op(N1799_t1) );
fim FAN_N1799_2 ( .fault(fault), .net(N1799), .FEN(FEN[767]), .op(N1799_t2) );
fim FAN_N1799_3 ( .fault(fault), .net(N1799), .FEN(FEN[768]), .op(N1799_t3) );
fim FAN_N1799_4 ( .fault(fault), .net(N1799), .FEN(FEN[769]), .op(N1799_t4) );
fim FAN_N1805_0 ( .fault(fault), .net(N1805), .FEN(FEN[770]), .op(N1805_t0) );
fim FAN_N1805_1 ( .fault(fault), .net(N1805), .FEN(FEN[771]), .op(N1805_t1) );
fim FAN_N1805_2 ( .fault(fault), .net(N1805), .FEN(FEN[772]), .op(N1805_t2) );
fim FAN_N1805_3 ( .fault(fault), .net(N1805), .FEN(FEN[773]), .op(N1805_t3) );
fim FAN_N1805_4 ( .fault(fault), .net(N1805), .FEN(FEN[774]), .op(N1805_t4) );
fim FAN_N2074_0 ( .fault(fault), .net(N2074), .FEN(FEN[775]), .op(N2074_t0) );
fim FAN_N2074_1 ( .fault(fault), .net(N2074), .FEN(FEN[776]), .op(N2074_t1) );
fim FAN_N2081_0 ( .fault(fault), .net(N2081), .FEN(FEN[777]), .op(N2081_t0) );
fim FAN_N2081_1 ( .fault(fault), .net(N2081), .FEN(FEN[778]), .op(N2081_t1) );
fim FAN_N141_0 ( .fault(fault), .net(N141), .FEN(FEN[779]), .op(N141_t0) );
fim FAN_N141_1 ( .fault(fault), .net(N141), .FEN(FEN[780]), .op(N141_t1) );
fim FAN_N1845_0 ( .fault(fault), .net(N1845), .FEN(FEN[781]), .op(N1845_t0) );
fim FAN_N1845_1 ( .fault(fault), .net(N1845), .FEN(FEN[782]), .op(N1845_t1) );
fim FAN_N1845_2 ( .fault(fault), .net(N1845), .FEN(FEN[783]), .op(N1845_t2) );
fim FAN_N1845_3 ( .fault(fault), .net(N1845), .FEN(FEN[784]), .op(N1845_t3) );
fim FAN_N1845_4 ( .fault(fault), .net(N1845), .FEN(FEN[785]), .op(N1845_t4) );
fim FAN_N147_0 ( .fault(fault), .net(N147), .FEN(FEN[786]), .op(N147_t0) );
fim FAN_N147_1 ( .fault(fault), .net(N147), .FEN(FEN[787]), .op(N147_t1) );
fim FAN_N138_0 ( .fault(fault), .net(N138), .FEN(FEN[788]), .op(N138_t0) );
fim FAN_N138_1 ( .fault(fault), .net(N138), .FEN(FEN[789]), .op(N138_t1) );
fim FAN_N144_0 ( .fault(fault), .net(N144), .FEN(FEN[790]), .op(N144_t0) );
fim FAN_N144_1 ( .fault(fault), .net(N144), .FEN(FEN[791]), .op(N144_t1) );
fim FAN_N135_0 ( .fault(fault), .net(N135), .FEN(FEN[792]), .op(N135_t0) );
fim FAN_N135_1 ( .fault(fault), .net(N135), .FEN(FEN[793]), .op(N135_t1) );
fim FAN_N1851_0 ( .fault(fault), .net(N1851), .FEN(FEN[794]), .op(N1851_t0) );
fim FAN_N1851_1 ( .fault(fault), .net(N1851), .FEN(FEN[795]), .op(N1851_t1) );
fim FAN_N1851_2 ( .fault(fault), .net(N1851), .FEN(FEN[796]), .op(N1851_t2) );
fim FAN_N1851_3 ( .fault(fault), .net(N1851), .FEN(FEN[797]), .op(N1851_t3) );
fim FAN_N1851_4 ( .fault(fault), .net(N1851), .FEN(FEN[798]), .op(N1851_t4) );
fim FAN_N1885_0 ( .fault(fault), .net(N1885), .FEN(FEN[799]), .op(N1885_t0) );
fim FAN_N1885_1 ( .fault(fault), .net(N1885), .FEN(FEN[800]), .op(N1885_t1) );
fim FAN_N1885_2 ( .fault(fault), .net(N1885), .FEN(FEN[801]), .op(N1885_t2) );
fim FAN_N1885_3 ( .fault(fault), .net(N1885), .FEN(FEN[802]), .op(N1885_t3) );
fim FAN_N1885_4 ( .fault(fault), .net(N1885), .FEN(FEN[803]), .op(N1885_t4) );
fim FAN_N1885_5 ( .fault(fault), .net(N1885), .FEN(FEN[804]), .op(N1885_t5) );
fim FAN_N1892_0 ( .fault(fault), .net(N1892), .FEN(FEN[805]), .op(N1892_t0) );
fim FAN_N1892_1 ( .fault(fault), .net(N1892), .FEN(FEN[806]), .op(N1892_t1) );
fim FAN_N1892_2 ( .fault(fault), .net(N1892), .FEN(FEN[807]), .op(N1892_t2) );
fim FAN_N1892_3 ( .fault(fault), .net(N1892), .FEN(FEN[808]), .op(N1892_t3) );
fim FAN_N1892_4 ( .fault(fault), .net(N1892), .FEN(FEN[809]), .op(N1892_t4) );
fim FAN_N1892_5 ( .fault(fault), .net(N1892), .FEN(FEN[810]), .op(N1892_t5) );
fim FAN_N103_0 ( .fault(fault), .net(N103), .FEN(FEN[811]), .op(N103_t0) );
fim FAN_N103_1 ( .fault(fault), .net(N103), .FEN(FEN[812]), .op(N103_t1) );
fim FAN_N130_0 ( .fault(fault), .net(N130), .FEN(FEN[813]), .op(N130_t0) );
fim FAN_N130_1 ( .fault(fault), .net(N130), .FEN(FEN[814]), .op(N130_t1) );
fim FAN_N127_0 ( .fault(fault), .net(N127), .FEN(FEN[815]), .op(N127_t0) );
fim FAN_N127_1 ( .fault(fault), .net(N127), .FEN(FEN[816]), .op(N127_t1) );
fim FAN_N124_0 ( .fault(fault), .net(N124), .FEN(FEN[817]), .op(N124_t0) );
fim FAN_N124_1 ( .fault(fault), .net(N124), .FEN(FEN[818]), .op(N124_t1) );
fim FAN_N100_0 ( .fault(fault), .net(N100), .FEN(FEN[819]), .op(N100_t0) );
fim FAN_N100_1 ( .fault(fault), .net(N100), .FEN(FEN[820]), .op(N100_t1) );
fim FAN_N1899_0 ( .fault(fault), .net(N1899), .FEN(FEN[821]), .op(N1899_t0) );
fim FAN_N1899_1 ( .fault(fault), .net(N1899), .FEN(FEN[822]), .op(N1899_t1) );
fim FAN_N1899_2 ( .fault(fault), .net(N1899), .FEN(FEN[823]), .op(N1899_t2) );
fim FAN_N1899_3 ( .fault(fault), .net(N1899), .FEN(FEN[824]), .op(N1899_t3) );
fim FAN_N1899_4 ( .fault(fault), .net(N1899), .FEN(FEN[825]), .op(N1899_t4) );
fim FAN_N1899_5 ( .fault(fault), .net(N1899), .FEN(FEN[826]), .op(N1899_t5) );
fim FAN_N1906_0 ( .fault(fault), .net(N1906), .FEN(FEN[827]), .op(N1906_t0) );
fim FAN_N1906_1 ( .fault(fault), .net(N1906), .FEN(FEN[828]), .op(N1906_t1) );
fim FAN_N1906_2 ( .fault(fault), .net(N1906), .FEN(FEN[829]), .op(N1906_t2) );
fim FAN_N1906_3 ( .fault(fault), .net(N1906), .FEN(FEN[830]), .op(N1906_t3) );
fim FAN_N1906_4 ( .fault(fault), .net(N1906), .FEN(FEN[831]), .op(N1906_t4) );
fim FAN_N1906_5 ( .fault(fault), .net(N1906), .FEN(FEN[832]), .op(N1906_t5) );
fim FAN_N115_0 ( .fault(fault), .net(N115), .FEN(FEN[833]), .op(N115_t0) );
fim FAN_N115_1 ( .fault(fault), .net(N115), .FEN(FEN[834]), .op(N115_t1) );
fim FAN_N118_0 ( .fault(fault), .net(N118), .FEN(FEN[835]), .op(N118_t0) );
fim FAN_N118_1 ( .fault(fault), .net(N118), .FEN(FEN[836]), .op(N118_t1) );
fim FAN_N97_0 ( .fault(fault), .net(N97), .FEN(FEN[837]), .op(N97_t0) );
fim FAN_N97_1 ( .fault(fault), .net(N97), .FEN(FEN[838]), .op(N97_t1) );
fim FAN_N94_0 ( .fault(fault), .net(N94), .FEN(FEN[839]), .op(N94_t0) );
fim FAN_N94_1 ( .fault(fault), .net(N94), .FEN(FEN[840]), .op(N94_t1) );
fim FAN_N121_0 ( .fault(fault), .net(N121), .FEN(FEN[841]), .op(N121_t0) );
fim FAN_N121_1 ( .fault(fault), .net(N121), .FEN(FEN[842]), .op(N121_t1) );
fim FAN_N1919_0 ( .fault(fault), .net(N1919), .FEN(FEN[843]), .op(N1919_t0) );
fim FAN_N1919_1 ( .fault(fault), .net(N1919), .FEN(FEN[844]), .op(N1919_t1) );
fim FAN_N1919_2 ( .fault(fault), .net(N1919), .FEN(FEN[845]), .op(N1919_t2) );
fim FAN_N1919_3 ( .fault(fault), .net(N1919), .FEN(FEN[846]), .op(N1919_t3) );
fim FAN_N1919_4 ( .fault(fault), .net(N1919), .FEN(FEN[847]), .op(N1919_t4) );
fim FAN_N1919_5 ( .fault(fault), .net(N1919), .FEN(FEN[848]), .op(N1919_t5) );
fim FAN_N1913_0 ( .fault(fault), .net(N1913), .FEN(FEN[849]), .op(N1913_t0) );
fim FAN_N1913_1 ( .fault(fault), .net(N1913), .FEN(FEN[850]), .op(N1913_t1) );
fim FAN_N1913_2 ( .fault(fault), .net(N1913), .FEN(FEN[851]), .op(N1913_t2) );
fim FAN_N1913_3 ( .fault(fault), .net(N1913), .FEN(FEN[852]), .op(N1913_t3) );
fim FAN_N1913_4 ( .fault(fault), .net(N1913), .FEN(FEN[853]), .op(N1913_t4) );
fim FAN_N1947_0 ( .fault(fault), .net(N1947), .FEN(FEN[854]), .op(N1947_t0) );
fim FAN_N1947_1 ( .fault(fault), .net(N1947), .FEN(FEN[855]), .op(N1947_t1) );
fim FAN_N1947_2 ( .fault(fault), .net(N1947), .FEN(FEN[856]), .op(N1947_t2) );
fim FAN_N1947_3 ( .fault(fault), .net(N1947), .FEN(FEN[857]), .op(N1947_t3) );
fim FAN_N1947_4 ( .fault(fault), .net(N1947), .FEN(FEN[858]), .op(N1947_t4) );
fim FAN_N1953_0 ( .fault(fault), .net(N1953), .FEN(FEN[859]), .op(N1953_t0) );
fim FAN_N1953_1 ( .fault(fault), .net(N1953), .FEN(FEN[860]), .op(N1953_t1) );
fim FAN_N1953_2 ( .fault(fault), .net(N1953), .FEN(FEN[861]), .op(N1953_t2) );
fim FAN_N2086_0 ( .fault(fault), .net(N2086), .FEN(FEN[862]), .op(N2086_t0) );
fim FAN_N2086_1 ( .fault(fault), .net(N2086), .FEN(FEN[863]), .op(N2086_t1) );
fim FAN_N1977_0 ( .fault(fault), .net(N1977), .FEN(FEN[864]), .op(N1977_t0) );
fim FAN_N1977_1 ( .fault(fault), .net(N1977), .FEN(FEN[865]), .op(N1977_t1) );
fim FAN_N1977_2 ( .fault(fault), .net(N1977), .FEN(FEN[866]), .op(N1977_t2) );
fim FAN_N1977_3 ( .fault(fault), .net(N1977), .FEN(FEN[867]), .op(N1977_t3) );
fim FAN_N1977_4 ( .fault(fault), .net(N1977), .FEN(FEN[868]), .op(N1977_t4) );
fim FAN_N1983_0 ( .fault(fault), .net(N1983), .FEN(FEN[869]), .op(N1983_t0) );
fim FAN_N1983_1 ( .fault(fault), .net(N1983), .FEN(FEN[870]), .op(N1983_t1) );
fim FAN_N1983_2 ( .fault(fault), .net(N1983), .FEN(FEN[871]), .op(N1983_t2) );
fim FAN_N1983_3 ( .fault(fault), .net(N1983), .FEN(FEN[872]), .op(N1983_t3) );
fim FAN_N1983_4 ( .fault(fault), .net(N1983), .FEN(FEN[873]), .op(N1983_t4) );
fim FAN_N759_0 ( .fault(fault), .net(N759), .FEN(FEN[874]), .op(N759_t0) );
fim FAN_N759_1 ( .fault(fault), .net(N759), .FEN(FEN[875]), .op(N759_t1) );
fim FAN_N70_0 ( .fault(fault), .net(N70), .FEN(FEN[876]), .op(N70_t0) );
fim FAN_N70_1 ( .fault(fault), .net(N70), .FEN(FEN[877]), .op(N70_t1) );
fim FAN_N2003_0 ( .fault(fault), .net(N2003), .FEN(FEN[878]), .op(N2003_t0) );
fim FAN_N2003_1 ( .fault(fault), .net(N2003), .FEN(FEN[879]), .op(N2003_t1) );
fim FAN_N2003_2 ( .fault(fault), .net(N2003), .FEN(FEN[880]), .op(N2003_t2) );
fim FAN_N2003_3 ( .fault(fault), .net(N2003), .FEN(FEN[881]), .op(N2003_t3) );
fim FAN_N2003_4 ( .fault(fault), .net(N2003), .FEN(FEN[882]), .op(N2003_t4) );
fim FAN_N2003_5 ( .fault(fault), .net(N2003), .FEN(FEN[883]), .op(N2003_t5) );
fim FAN_N1997_0 ( .fault(fault), .net(N1997), .FEN(FEN[884]), .op(N1997_t0) );
fim FAN_N1997_1 ( .fault(fault), .net(N1997), .FEN(FEN[885]), .op(N1997_t1) );
fim FAN_N1997_2 ( .fault(fault), .net(N1997), .FEN(FEN[886]), .op(N1997_t2) );
fim FAN_N1997_3 ( .fault(fault), .net(N1997), .FEN(FEN[887]), .op(N1997_t3) );
fim FAN_N1997_4 ( .fault(fault), .net(N1997), .FEN(FEN[888]), .op(N1997_t4) );
fim FAN_N2024_0 ( .fault(fault), .net(N2024), .FEN(FEN[889]), .op(N2024_t0) );
fim FAN_N2024_1 ( .fault(fault), .net(N2024), .FEN(FEN[890]), .op(N2024_t1) );
fim FAN_N2024_2 ( .fault(fault), .net(N2024), .FEN(FEN[891]), .op(N2024_t2) );
fim FAN_N2024_3 ( .fault(fault), .net(N2024), .FEN(FEN[892]), .op(N2024_t3) );
fim FAN_N2024_4 ( .fault(fault), .net(N2024), .FEN(FEN[893]), .op(N2024_t4) );
fim FAN_N2024_5 ( .fault(fault), .net(N2024), .FEN(FEN[894]), .op(N2024_t5) );
fim FAN_N2031_0 ( .fault(fault), .net(N2031), .FEN(FEN[895]), .op(N2031_t0) );
fim FAN_N2031_1 ( .fault(fault), .net(N2031), .FEN(FEN[896]), .op(N2031_t1) );
fim FAN_N2031_2 ( .fault(fault), .net(N2031), .FEN(FEN[897]), .op(N2031_t2) );
fim FAN_N2031_3 ( .fault(fault), .net(N2031), .FEN(FEN[898]), .op(N2031_t3) );
fim FAN_N2031_4 ( .fault(fault), .net(N2031), .FEN(FEN[899]), .op(N2031_t4) );
fim FAN_N2031_5 ( .fault(fault), .net(N2031), .FEN(FEN[900]), .op(N2031_t5) );
fim FAN_N2038_0 ( .fault(fault), .net(N2038), .FEN(FEN[901]), .op(N2038_t0) );
fim FAN_N2038_1 ( .fault(fault), .net(N2038), .FEN(FEN[902]), .op(N2038_t1) );
fim FAN_N2038_2 ( .fault(fault), .net(N2038), .FEN(FEN[903]), .op(N2038_t2) );
fim FAN_N2038_3 ( .fault(fault), .net(N2038), .FEN(FEN[904]), .op(N2038_t3) );
fim FAN_N2038_4 ( .fault(fault), .net(N2038), .FEN(FEN[905]), .op(N2038_t4) );
fim FAN_N2038_5 ( .fault(fault), .net(N2038), .FEN(FEN[906]), .op(N2038_t5) );
fim FAN_N2045_0 ( .fault(fault), .net(N2045), .FEN(FEN[907]), .op(N2045_t0) );
fim FAN_N2045_1 ( .fault(fault), .net(N2045), .FEN(FEN[908]), .op(N2045_t1) );
fim FAN_N2045_2 ( .fault(fault), .net(N2045), .FEN(FEN[909]), .op(N2045_t2) );
fim FAN_N2045_3 ( .fault(fault), .net(N2045), .FEN(FEN[910]), .op(N2045_t3) );
fim FAN_N2045_4 ( .fault(fault), .net(N2045), .FEN(FEN[911]), .op(N2045_t4) );
fim FAN_N2045_5 ( .fault(fault), .net(N2045), .FEN(FEN[912]), .op(N2045_t5) );
fim FAN_N2052_0 ( .fault(fault), .net(N2052), .FEN(FEN[913]), .op(N2052_t0) );
fim FAN_N2052_1 ( .fault(fault), .net(N2052), .FEN(FEN[914]), .op(N2052_t1) );
fim FAN_N2052_2 ( .fault(fault), .net(N2052), .FEN(FEN[915]), .op(N2052_t2) );
fim FAN_N2052_3 ( .fault(fault), .net(N2052), .FEN(FEN[916]), .op(N2052_t3) );
fim FAN_N2052_4 ( .fault(fault), .net(N2052), .FEN(FEN[917]), .op(N2052_t4) );
fim FAN_N2058_0 ( .fault(fault), .net(N2058), .FEN(FEN[918]), .op(N2058_t0) );
fim FAN_N2058_1 ( .fault(fault), .net(N2058), .FEN(FEN[919]), .op(N2058_t1) );
fim FAN_N2058_2 ( .fault(fault), .net(N2058), .FEN(FEN[920]), .op(N2058_t2) );
fim FAN_N2058_3 ( .fault(fault), .net(N2058), .FEN(FEN[921]), .op(N2058_t3) );
fim FAN_N2058_4 ( .fault(fault), .net(N2058), .FEN(FEN[922]), .op(N2058_t4) );
fim FAN_N1119_0 ( .fault(fault), .net(N1119), .FEN(FEN[923]), .op(N1119_t0) );
fim FAN_N1119_1 ( .fault(fault), .net(N1119), .FEN(FEN[924]), .op(N1119_t1) );
fim FAN_N1119_2 ( .fault(fault), .net(N1119), .FEN(FEN[925]), .op(N1119_t2) );
fim FAN_N1119_3 ( .fault(fault), .net(N1119), .FEN(FEN[926]), .op(N1119_t3) );
fim FAN_N1119_4 ( .fault(fault), .net(N1119), .FEN(FEN[927]), .op(N1119_t4) );
fim FAN_N1132_0 ( .fault(fault), .net(N1132), .FEN(FEN[928]), .op(N1132_t0) );
fim FAN_N1132_1 ( .fault(fault), .net(N1132), .FEN(FEN[929]), .op(N1132_t1) );
fim FAN_N1132_2 ( .fault(fault), .net(N1132), .FEN(FEN[930]), .op(N1132_t2) );
fim FAN_N1141_0 ( .fault(fault), .net(N1141), .FEN(FEN[931]), .op(N1141_t0) );
fim FAN_N1141_1 ( .fault(fault), .net(N1141), .FEN(FEN[932]), .op(N1141_t1) );
fim FAN_N1141_2 ( .fault(fault), .net(N1141), .FEN(FEN[933]), .op(N1141_t2) );
fim FAN_N1141_3 ( .fault(fault), .net(N1141), .FEN(FEN[934]), .op(N1141_t3) );
fim FAN_N1141_4 ( .fault(fault), .net(N1141), .FEN(FEN[935]), .op(N1141_t4) );
fim FAN_N1154_0 ( .fault(fault), .net(N1154), .FEN(FEN[936]), .op(N1154_t0) );
fim FAN_N1154_1 ( .fault(fault), .net(N1154), .FEN(FEN[937]), .op(N1154_t1) );
fim FAN_N1154_2 ( .fault(fault), .net(N1154), .FEN(FEN[938]), .op(N1154_t2) );
fim FAN_N1154_3 ( .fault(fault), .net(N1154), .FEN(FEN[939]), .op(N1154_t3) );
fim FAN_N1154_4 ( .fault(fault), .net(N1154), .FEN(FEN[940]), .op(N1154_t4) );
fim FAN_N2235_0 ( .fault(fault), .net(N2235), .FEN(FEN[941]), .op(N2235_t0) );
fim FAN_N2235_1 ( .fault(fault), .net(N2235), .FEN(FEN[942]), .op(N2235_t1) );
fim FAN_N1227_0 ( .fault(fault), .net(N1227), .FEN(FEN[943]), .op(N1227_t0) );
fim FAN_N1227_1 ( .fault(fault), .net(N1227), .FEN(FEN[944]), .op(N1227_t1) );
fim FAN_N1227_2 ( .fault(fault), .net(N1227), .FEN(FEN[945]), .op(N1227_t2) );
fim FAN_N1227_3 ( .fault(fault), .net(N1227), .FEN(FEN[946]), .op(N1227_t3) );
fim FAN_N1227_4 ( .fault(fault), .net(N1227), .FEN(FEN[947]), .op(N1227_t4) );
fim FAN_N1240_0 ( .fault(fault), .net(N1240), .FEN(FEN[948]), .op(N1240_t0) );
fim FAN_N1240_1 ( .fault(fault), .net(N1240), .FEN(FEN[949]), .op(N1240_t1) );
fim FAN_N1240_2 ( .fault(fault), .net(N1240), .FEN(FEN[950]), .op(N1240_t2) );
fim FAN_N2231_0 ( .fault(fault), .net(N2231), .FEN(FEN[951]), .op(N2231_t0) );
fim FAN_N2231_1 ( .fault(fault), .net(N2231), .FEN(FEN[952]), .op(N2231_t1) );
fim FAN_N2257_0 ( .fault(fault), .net(N2257), .FEN(FEN[953]), .op(N2257_t0) );
fim FAN_N2257_1 ( .fault(fault), .net(N2257), .FEN(FEN[954]), .op(N2257_t1) );
fim FAN_N2257_2 ( .fault(fault), .net(N2257), .FEN(FEN[955]), .op(N2257_t2) );
fim FAN_N2257_3 ( .fault(fault), .net(N2257), .FEN(FEN[956]), .op(N2257_t3) );
fim FAN_N2257_4 ( .fault(fault), .net(N2257), .FEN(FEN[957]), .op(N2257_t4) );
fim FAN_N2257_5 ( .fault(fault), .net(N2257), .FEN(FEN[958]), .op(N2257_t5) );
fim FAN_N2257_6 ( .fault(fault), .net(N2257), .FEN(FEN[959]), .op(N2257_t6) );
fim FAN_N2257_7 ( .fault(fault), .net(N2257), .FEN(FEN[960]), .op(N2257_t7) );
fim FAN_N2257_8 ( .fault(fault), .net(N2257), .FEN(FEN[961]), .op(N2257_t8) );
fim FAN_N2269_0 ( .fault(fault), .net(N2269), .FEN(FEN[962]), .op(N2269_t0) );
fim FAN_N2269_1 ( .fault(fault), .net(N2269), .FEN(FEN[963]), .op(N2269_t1) );
fim FAN_N2269_2 ( .fault(fault), .net(N2269), .FEN(FEN[964]), .op(N2269_t2) );
fim FAN_N2269_3 ( .fault(fault), .net(N2269), .FEN(FEN[965]), .op(N2269_t3) );
fim FAN_N2287_0 ( .fault(fault), .net(N2287), .FEN(FEN[966]), .op(N2287_t0) );
fim FAN_N2287_1 ( .fault(fault), .net(N2287), .FEN(FEN[967]), .op(N2287_t1) );
fim FAN_N2287_2 ( .fault(fault), .net(N2287), .FEN(FEN[968]), .op(N2287_t2) );
fim FAN_N2287_3 ( .fault(fault), .net(N2287), .FEN(FEN[969]), .op(N2287_t3) );
fim FAN_N2287_4 ( .fault(fault), .net(N2287), .FEN(FEN[970]), .op(N2287_t4) );
fim FAN_N2293_0 ( .fault(fault), .net(N2293), .FEN(FEN[971]), .op(N2293_t0) );
fim FAN_N2293_1 ( .fault(fault), .net(N2293), .FEN(FEN[972]), .op(N2293_t1) );
fim FAN_N2293_2 ( .fault(fault), .net(N2293), .FEN(FEN[973]), .op(N2293_t2) );
fim FAN_N2293_3 ( .fault(fault), .net(N2293), .FEN(FEN[974]), .op(N2293_t3) );
fim FAN_N2293_4 ( .fault(fault), .net(N2293), .FEN(FEN[975]), .op(N2293_t4) );
fim FAN_N2309_0 ( .fault(fault), .net(N2309), .FEN(FEN[976]), .op(N2309_t0) );
fim FAN_N2309_1 ( .fault(fault), .net(N2309), .FEN(FEN[977]), .op(N2309_t1) );
fim FAN_N2309_2 ( .fault(fault), .net(N2309), .FEN(FEN[978]), .op(N2309_t2) );
fim FAN_N2309_3 ( .fault(fault), .net(N2309), .FEN(FEN[979]), .op(N2309_t3) );
fim FAN_N2309_4 ( .fault(fault), .net(N2309), .FEN(FEN[980]), .op(N2309_t4) );
fim FAN_N2315_0 ( .fault(fault), .net(N2315), .FEN(FEN[981]), .op(N2315_t0) );
fim FAN_N2315_1 ( .fault(fault), .net(N2315), .FEN(FEN[982]), .op(N2315_t1) );
fim FAN_N2315_2 ( .fault(fault), .net(N2315), .FEN(FEN[983]), .op(N2315_t2) );
fim FAN_N2315_3 ( .fault(fault), .net(N2315), .FEN(FEN[984]), .op(N2315_t3) );
fim FAN_N2315_4 ( .fault(fault), .net(N2315), .FEN(FEN[985]), .op(N2315_t4) );
fim FAN_N2331_0 ( .fault(fault), .net(N2331), .FEN(FEN[986]), .op(N2331_t0) );
fim FAN_N2331_1 ( .fault(fault), .net(N2331), .FEN(FEN[987]), .op(N2331_t1) );
fim FAN_N2331_2 ( .fault(fault), .net(N2331), .FEN(FEN[988]), .op(N2331_t2) );
fim FAN_N2331_3 ( .fault(fault), .net(N2331), .FEN(FEN[989]), .op(N2331_t3) );
fim FAN_N2331_4 ( .fault(fault), .net(N2331), .FEN(FEN[990]), .op(N2331_t4) );
fim FAN_N2368_0 ( .fault(fault), .net(N2368), .FEN(FEN[991]), .op(N2368_t0) );
fim FAN_N2368_1 ( .fault(fault), .net(N2368), .FEN(FEN[992]), .op(N2368_t1) );
fim FAN_N2368_2 ( .fault(fault), .net(N2368), .FEN(FEN[993]), .op(N2368_t2) );
fim FAN_N2368_3 ( .fault(fault), .net(N2368), .FEN(FEN[994]), .op(N2368_t3) );
fim FAN_N2368_4 ( .fault(fault), .net(N2368), .FEN(FEN[995]), .op(N2368_t4) );
fim FAN_N2384_0 ( .fault(fault), .net(N2384), .FEN(FEN[996]), .op(N2384_t0) );
fim FAN_N2384_1 ( .fault(fault), .net(N2384), .FEN(FEN[997]), .op(N2384_t1) );
fim FAN_N2384_2 ( .fault(fault), .net(N2384), .FEN(FEN[998]), .op(N2384_t2) );
fim FAN_N2384_3 ( .fault(fault), .net(N2384), .FEN(FEN[999]), .op(N2384_t3) );
fim FAN_N2384_4 ( .fault(fault), .net(N2384), .FEN(FEN[1000]), .op(N2384_t4) );
fim FAN_N2390_0 ( .fault(fault), .net(N2390), .FEN(FEN[1001]), .op(N2390_t0) );
fim FAN_N2390_1 ( .fault(fault), .net(N2390), .FEN(FEN[1002]), .op(N2390_t1) );
fim FAN_N2390_2 ( .fault(fault), .net(N2390), .FEN(FEN[1003]), .op(N2390_t2) );
fim FAN_N2390_3 ( .fault(fault), .net(N2390), .FEN(FEN[1004]), .op(N2390_t3) );
fim FAN_N2390_4 ( .fault(fault), .net(N2390), .FEN(FEN[1005]), .op(N2390_t4) );
fim FAN_N2406_0 ( .fault(fault), .net(N2406), .FEN(FEN[1006]), .op(N2406_t0) );
fim FAN_N2406_1 ( .fault(fault), .net(N2406), .FEN(FEN[1007]), .op(N2406_t1) );
fim FAN_N2406_2 ( .fault(fault), .net(N2406), .FEN(FEN[1008]), .op(N2406_t2) );
fim FAN_N2406_3 ( .fault(fault), .net(N2406), .FEN(FEN[1009]), .op(N2406_t3) );
fim FAN_N2406_4 ( .fault(fault), .net(N2406), .FEN(FEN[1010]), .op(N2406_t4) );
fim FAN_N2412_0 ( .fault(fault), .net(N2412), .FEN(FEN[1011]), .op(N2412_t0) );
fim FAN_N2412_1 ( .fault(fault), .net(N2412), .FEN(FEN[1012]), .op(N2412_t1) );
fim FAN_N2412_2 ( .fault(fault), .net(N2412), .FEN(FEN[1013]), .op(N2412_t2) );
fim FAN_N2412_3 ( .fault(fault), .net(N2412), .FEN(FEN[1014]), .op(N2412_t3) );
fim FAN_N2412_4 ( .fault(fault), .net(N2412), .FEN(FEN[1015]), .op(N2412_t4) );
fim FAN_N2644_0 ( .fault(fault), .net(N2644), .FEN(FEN[1016]), .op(N2644_t0) );
fim FAN_N2644_1 ( .fault(fault), .net(N2644), .FEN(FEN[1017]), .op(N2644_t1) );
fim FAN_N2644_2 ( .fault(fault), .net(N2644), .FEN(FEN[1018]), .op(N2644_t2) );
fim FAN_N2644_3 ( .fault(fault), .net(N2644), .FEN(FEN[1019]), .op(N2644_t3) );
fim FAN_N2644_4 ( .fault(fault), .net(N2644), .FEN(FEN[1020]), .op(N2644_t4) );
fim FAN_N2638_0 ( .fault(fault), .net(N2638), .FEN(FEN[1021]), .op(N2638_t0) );
fim FAN_N2638_1 ( .fault(fault), .net(N2638), .FEN(FEN[1022]), .op(N2638_t1) );
fim FAN_N2638_2 ( .fault(fault), .net(N2638), .FEN(FEN[1023]), .op(N2638_t2) );
fim FAN_N2638_3 ( .fault(fault), .net(N2638), .FEN(FEN[1024]), .op(N2638_t3) );
fim FAN_N2638_4 ( .fault(fault), .net(N2638), .FEN(FEN[1025]), .op(N2638_t4) );
fim FAN_N2632_0 ( .fault(fault), .net(N2632), .FEN(FEN[1026]), .op(N2632_t0) );
fim FAN_N2632_1 ( .fault(fault), .net(N2632), .FEN(FEN[1027]), .op(N2632_t1) );
fim FAN_N2632_2 ( .fault(fault), .net(N2632), .FEN(FEN[1028]), .op(N2632_t2) );
fim FAN_N2632_3 ( .fault(fault), .net(N2632), .FEN(FEN[1029]), .op(N2632_t3) );
fim FAN_N2632_4 ( .fault(fault), .net(N2632), .FEN(FEN[1030]), .op(N2632_t4) );
fim FAN_N2626_0 ( .fault(fault), .net(N2626), .FEN(FEN[1031]), .op(N2626_t0) );
fim FAN_N2626_1 ( .fault(fault), .net(N2626), .FEN(FEN[1032]), .op(N2626_t1) );
fim FAN_N2626_2 ( .fault(fault), .net(N2626), .FEN(FEN[1033]), .op(N2626_t2) );
fim FAN_N2626_3 ( .fault(fault), .net(N2626), .FEN(FEN[1034]), .op(N2626_t3) );
fim FAN_N2626_4 ( .fault(fault), .net(N2626), .FEN(FEN[1035]), .op(N2626_t4) );
fim FAN_N2619_0 ( .fault(fault), .net(N2619), .FEN(FEN[1036]), .op(N2619_t0) );
fim FAN_N2619_1 ( .fault(fault), .net(N2619), .FEN(FEN[1037]), .op(N2619_t1) );
fim FAN_N2619_2 ( .fault(fault), .net(N2619), .FEN(FEN[1038]), .op(N2619_t2) );
fim FAN_N2619_3 ( .fault(fault), .net(N2619), .FEN(FEN[1039]), .op(N2619_t3) );
fim FAN_N2619_4 ( .fault(fault), .net(N2619), .FEN(FEN[1040]), .op(N2619_t4) );
fim FAN_N2619_5 ( .fault(fault), .net(N2619), .FEN(FEN[1041]), .op(N2619_t5) );
fim FAN_N2523_0 ( .fault(fault), .net(N2523), .FEN(FEN[1042]), .op(N2523_t0) );
fim FAN_N2523_1 ( .fault(fault), .net(N2523), .FEN(FEN[1043]), .op(N2523_t1) );
fim FAN_N2523_2 ( .fault(fault), .net(N2523), .FEN(FEN[1044]), .op(N2523_t2) );
fim FAN_N2523_3 ( .fault(fault), .net(N2523), .FEN(FEN[1045]), .op(N2523_t3) );
fim FAN_N2523_4 ( .fault(fault), .net(N2523), .FEN(FEN[1046]), .op(N2523_t4) );
fim FAN_N1167_0 ( .fault(fault), .net(N1167), .FEN(FEN[1047]), .op(N1167_t0) );
fim FAN_N1167_1 ( .fault(fault), .net(N1167), .FEN(FEN[1048]), .op(N1167_t1) );
fim FAN_N1167_2 ( .fault(fault), .net(N1167), .FEN(FEN[1049]), .op(N1167_t2) );
fim FAN_N1167_3 ( .fault(fault), .net(N1167), .FEN(FEN[1050]), .op(N1167_t3) );
fim FAN_N2533_0 ( .fault(fault), .net(N2533), .FEN(FEN[1051]), .op(N2533_t0) );
fim FAN_N2533_1 ( .fault(fault), .net(N2533), .FEN(FEN[1052]), .op(N2533_t1) );
fim FAN_N2533_2 ( .fault(fault), .net(N2533), .FEN(FEN[1053]), .op(N2533_t2) );
fim FAN_N2778_0 ( .fault(fault), .net(N2778), .FEN(FEN[1054]), .op(N2778_t0) );
fim FAN_N2778_1 ( .fault(fault), .net(N2778), .FEN(FEN[1055]), .op(N2778_t1) );
fim FAN_N2508_0 ( .fault(fault), .net(N2508), .FEN(FEN[1056]), .op(N2508_t0) );
fim FAN_N2508_1 ( .fault(fault), .net(N2508), .FEN(FEN[1057]), .op(N2508_t1) );
fim FAN_N2508_2 ( .fault(fault), .net(N2508), .FEN(FEN[1058]), .op(N2508_t2) );
fim FAN_N2508_3 ( .fault(fault), .net(N2508), .FEN(FEN[1059]), .op(N2508_t3) );
fim FAN_N2508_4 ( .fault(fault), .net(N2508), .FEN(FEN[1060]), .op(N2508_t4) );
fim FAN_N2502_0 ( .fault(fault), .net(N2502), .FEN(FEN[1061]), .op(N2502_t0) );
fim FAN_N2502_1 ( .fault(fault), .net(N2502), .FEN(FEN[1062]), .op(N2502_t1) );
fim FAN_N2502_2 ( .fault(fault), .net(N2502), .FEN(FEN[1063]), .op(N2502_t2) );
fim FAN_N2502_3 ( .fault(fault), .net(N2502), .FEN(FEN[1064]), .op(N2502_t3) );
fim FAN_N2502_4 ( .fault(fault), .net(N2502), .FEN(FEN[1065]), .op(N2502_t4) );
fim FAN_N2496_0 ( .fault(fault), .net(N2496), .FEN(FEN[1066]), .op(N2496_t0) );
fim FAN_N2496_1 ( .fault(fault), .net(N2496), .FEN(FEN[1067]), .op(N2496_t1) );
fim FAN_N2496_2 ( .fault(fault), .net(N2496), .FEN(FEN[1068]), .op(N2496_t2) );
fim FAN_N2496_3 ( .fault(fault), .net(N2496), .FEN(FEN[1069]), .op(N2496_t3) );
fim FAN_N2496_4 ( .fault(fault), .net(N2496), .FEN(FEN[1070]), .op(N2496_t4) );
fim FAN_N2488_0 ( .fault(fault), .net(N2488), .FEN(FEN[1071]), .op(N2488_t0) );
fim FAN_N2488_1 ( .fault(fault), .net(N2488), .FEN(FEN[1072]), .op(N2488_t1) );
fim FAN_N2488_2 ( .fault(fault), .net(N2488), .FEN(FEN[1073]), .op(N2488_t2) );
fim FAN_N2488_3 ( .fault(fault), .net(N2488), .FEN(FEN[1074]), .op(N2488_t3) );
fim FAN_N2488_4 ( .fault(fault), .net(N2488), .FEN(FEN[1075]), .op(N2488_t4) );
fim FAN_N2488_5 ( .fault(fault), .net(N2488), .FEN(FEN[1076]), .op(N2488_t5) );
fim FAN_N2488_6 ( .fault(fault), .net(N2488), .FEN(FEN[1077]), .op(N2488_t6) );
fim FAN_N2482_0 ( .fault(fault), .net(N2482), .FEN(FEN[1078]), .op(N2482_t0) );
fim FAN_N2482_1 ( .fault(fault), .net(N2482), .FEN(FEN[1079]), .op(N2482_t1) );
fim FAN_N2482_2 ( .fault(fault), .net(N2482), .FEN(FEN[1080]), .op(N2482_t2) );
fim FAN_N2482_3 ( .fault(fault), .net(N2482), .FEN(FEN[1081]), .op(N2482_t3) );
fim FAN_N2482_4 ( .fault(fault), .net(N2482), .FEN(FEN[1082]), .op(N2482_t4) );
fim FAN_N2573_0 ( .fault(fault), .net(N2573), .FEN(FEN[1083]), .op(N2573_t0) );
fim FAN_N2573_1 ( .fault(fault), .net(N2573), .FEN(FEN[1084]), .op(N2573_t1) );
fim FAN_N2573_2 ( .fault(fault), .net(N2573), .FEN(FEN[1085]), .op(N2573_t2) );
fim FAN_N2573_3 ( .fault(fault), .net(N2573), .FEN(FEN[1086]), .op(N2573_t3) );
fim FAN_N2573_4 ( .fault(fault), .net(N2573), .FEN(FEN[1087]), .op(N2573_t4) );
fim FAN_N2567_0 ( .fault(fault), .net(N2567), .FEN(FEN[1088]), .op(N2567_t0) );
fim FAN_N2567_1 ( .fault(fault), .net(N2567), .FEN(FEN[1089]), .op(N2567_t1) );
fim FAN_N2567_2 ( .fault(fault), .net(N2567), .FEN(FEN[1090]), .op(N2567_t2) );
fim FAN_N2567_3 ( .fault(fault), .net(N2567), .FEN(FEN[1091]), .op(N2567_t3) );
fim FAN_N2567_4 ( .fault(fault), .net(N2567), .FEN(FEN[1092]), .op(N2567_t4) );
fim FAN_N2561_0 ( .fault(fault), .net(N2561), .FEN(FEN[1093]), .op(N2561_t0) );
fim FAN_N2561_1 ( .fault(fault), .net(N2561), .FEN(FEN[1094]), .op(N2561_t1) );
fim FAN_N2561_2 ( .fault(fault), .net(N2561), .FEN(FEN[1095]), .op(N2561_t2) );
fim FAN_N2561_3 ( .fault(fault), .net(N2561), .FEN(FEN[1096]), .op(N2561_t3) );
fim FAN_N2561_4 ( .fault(fault), .net(N2561), .FEN(FEN[1097]), .op(N2561_t4) );
fim FAN_N2554_0 ( .fault(fault), .net(N2554), .FEN(FEN[1098]), .op(N2554_t0) );
fim FAN_N2554_1 ( .fault(fault), .net(N2554), .FEN(FEN[1099]), .op(N2554_t1) );
fim FAN_N2554_2 ( .fault(fault), .net(N2554), .FEN(FEN[1100]), .op(N2554_t2) );
fim FAN_N2554_3 ( .fault(fault), .net(N2554), .FEN(FEN[1101]), .op(N2554_t3) );
fim FAN_N2554_4 ( .fault(fault), .net(N2554), .FEN(FEN[1102]), .op(N2554_t4) );
fim FAN_N2554_5 ( .fault(fault), .net(N2554), .FEN(FEN[1103]), .op(N2554_t5) );
fim FAN_N2761_0 ( .fault(fault), .net(N2761), .FEN(FEN[1104]), .op(N2761_t0) );
fim FAN_N2761_1 ( .fault(fault), .net(N2761), .FEN(FEN[1105]), .op(N2761_t1) );
fim FAN_N2761_2 ( .fault(fault), .net(N2761), .FEN(FEN[1106]), .op(N2761_t2) );
fim FAN_N2478_0 ( .fault(fault), .net(N2478), .FEN(FEN[1107]), .op(N2478_t0) );
fim FAN_N2478_1 ( .fault(fault), .net(N2478), .FEN(FEN[1108]), .op(N2478_t1) );
fim FAN_N2478_2 ( .fault(fault), .net(N2478), .FEN(FEN[1109]), .op(N2478_t2) );
fim FAN_N2757_0 ( .fault(fault), .net(N2757), .FEN(FEN[1110]), .op(N2757_t0) );
fim FAN_N2757_1 ( .fault(fault), .net(N2757), .FEN(FEN[1111]), .op(N2757_t1) );
fim FAN_N2757_2 ( .fault(fault), .net(N2757), .FEN(FEN[1112]), .op(N2757_t2) );
fim FAN_N2474_0 ( .fault(fault), .net(N2474), .FEN(FEN[1113]), .op(N2474_t0) );
fim FAN_N2474_1 ( .fault(fault), .net(N2474), .FEN(FEN[1114]), .op(N2474_t1) );
fim FAN_N2474_2 ( .fault(fault), .net(N2474), .FEN(FEN[1115]), .op(N2474_t2) );
fim FAN_N2753_0 ( .fault(fault), .net(N2753), .FEN(FEN[1116]), .op(N2753_t0) );
fim FAN_N2753_1 ( .fault(fault), .net(N2753), .FEN(FEN[1117]), .op(N2753_t1) );
fim FAN_N2753_2 ( .fault(fault), .net(N2753), .FEN(FEN[1118]), .op(N2753_t2) );
fim FAN_N2470_0 ( .fault(fault), .net(N2470), .FEN(FEN[1119]), .op(N2470_t0) );
fim FAN_N2470_1 ( .fault(fault), .net(N2470), .FEN(FEN[1120]), .op(N2470_t1) );
fim FAN_N2470_2 ( .fault(fault), .net(N2470), .FEN(FEN[1121]), .op(N2470_t2) );
fim FAN_N2749_0 ( .fault(fault), .net(N2749), .FEN(FEN[1122]), .op(N2749_t0) );
fim FAN_N2749_1 ( .fault(fault), .net(N2749), .FEN(FEN[1123]), .op(N2749_t1) );
fim FAN_N2749_2 ( .fault(fault), .net(N2749), .FEN(FEN[1124]), .op(N2749_t2) );
fim FAN_N2466_0 ( .fault(fault), .net(N2466), .FEN(FEN[1125]), .op(N2466_t0) );
fim FAN_N2466_1 ( .fault(fault), .net(N2466), .FEN(FEN[1126]), .op(N2466_t1) );
fim FAN_N2466_2 ( .fault(fault), .net(N2466), .FEN(FEN[1127]), .op(N2466_t2) );
fim FAN_N2745_0 ( .fault(fault), .net(N2745), .FEN(FEN[1128]), .op(N2745_t0) );
fim FAN_N2745_1 ( .fault(fault), .net(N2745), .FEN(FEN[1129]), .op(N2745_t1) );
fim FAN_N2745_2 ( .fault(fault), .net(N2745), .FEN(FEN[1130]), .op(N2745_t2) );
fim FAN_N2462_0 ( .fault(fault), .net(N2462), .FEN(FEN[1131]), .op(N2462_t0) );
fim FAN_N2462_1 ( .fault(fault), .net(N2462), .FEN(FEN[1132]), .op(N2462_t1) );
fim FAN_N2462_2 ( .fault(fault), .net(N2462), .FEN(FEN[1133]), .op(N2462_t2) );
fim FAN_N2741_0 ( .fault(fault), .net(N2741), .FEN(FEN[1134]), .op(N2741_t0) );
fim FAN_N2741_1 ( .fault(fault), .net(N2741), .FEN(FEN[1135]), .op(N2741_t1) );
fim FAN_N2741_2 ( .fault(fault), .net(N2741), .FEN(FEN[1136]), .op(N2741_t2) );
fim FAN_N2550_0 ( .fault(fault), .net(N2550), .FEN(FEN[1137]), .op(N2550_t0) );
fim FAN_N2550_1 ( .fault(fault), .net(N2550), .FEN(FEN[1138]), .op(N2550_t1) );
fim FAN_N2550_2 ( .fault(fault), .net(N2550), .FEN(FEN[1139]), .op(N2550_t2) );
fim FAN_N2737_0 ( .fault(fault), .net(N2737), .FEN(FEN[1140]), .op(N2737_t0) );
fim FAN_N2737_1 ( .fault(fault), .net(N2737), .FEN(FEN[1141]), .op(N2737_t1) );
fim FAN_N2737_2 ( .fault(fault), .net(N2737), .FEN(FEN[1142]), .op(N2737_t2) );
fim FAN_N2546_0 ( .fault(fault), .net(N2546), .FEN(FEN[1143]), .op(N2546_t0) );
fim FAN_N2546_1 ( .fault(fault), .net(N2546), .FEN(FEN[1144]), .op(N2546_t1) );
fim FAN_N2546_2 ( .fault(fault), .net(N2546), .FEN(FEN[1145]), .op(N2546_t2) );
fim FAN_N2733_0 ( .fault(fault), .net(N2733), .FEN(FEN[1146]), .op(N2733_t0) );
fim FAN_N2733_1 ( .fault(fault), .net(N2733), .FEN(FEN[1147]), .op(N2733_t1) );
fim FAN_N2733_2 ( .fault(fault), .net(N2733), .FEN(FEN[1148]), .op(N2733_t2) );
fim FAN_N2542_0 ( .fault(fault), .net(N2542), .FEN(FEN[1149]), .op(N2542_t0) );
fim FAN_N2542_1 ( .fault(fault), .net(N2542), .FEN(FEN[1150]), .op(N2542_t1) );
fim FAN_N2542_2 ( .fault(fault), .net(N2542), .FEN(FEN[1151]), .op(N2542_t2) );
fim FAN_N2729_0 ( .fault(fault), .net(N2729), .FEN(FEN[1152]), .op(N2729_t0) );
fim FAN_N2729_1 ( .fault(fault), .net(N2729), .FEN(FEN[1153]), .op(N2729_t1) );
fim FAN_N2729_2 ( .fault(fault), .net(N2729), .FEN(FEN[1154]), .op(N2729_t2) );
fim FAN_N2538_0 ( .fault(fault), .net(N2538), .FEN(FEN[1155]), .op(N2538_t0) );
fim FAN_N2538_1 ( .fault(fault), .net(N2538), .FEN(FEN[1156]), .op(N2538_t1) );
fim FAN_N2538_2 ( .fault(fault), .net(N2538), .FEN(FEN[1157]), .op(N2538_t2) );
fim FAN_N2670_0 ( .fault(fault), .net(N2670), .FEN(FEN[1158]), .op(N2670_t0) );
fim FAN_N2670_1 ( .fault(fault), .net(N2670), .FEN(FEN[1159]), .op(N2670_t1) );
fim FAN_N2670_2 ( .fault(fault), .net(N2670), .FEN(FEN[1160]), .op(N2670_t2) );
fim FAN_N2458_0 ( .fault(fault), .net(N2458), .FEN(FEN[1161]), .op(N2458_t0) );
fim FAN_N2458_1 ( .fault(fault), .net(N2458), .FEN(FEN[1162]), .op(N2458_t1) );
fim FAN_N2458_2 ( .fault(fault), .net(N2458), .FEN(FEN[1163]), .op(N2458_t2) );
fim FAN_N2666_0 ( .fault(fault), .net(N2666), .FEN(FEN[1164]), .op(N2666_t0) );
fim FAN_N2666_1 ( .fault(fault), .net(N2666), .FEN(FEN[1165]), .op(N2666_t1) );
fim FAN_N2666_2 ( .fault(fault), .net(N2666), .FEN(FEN[1166]), .op(N2666_t2) );
fim FAN_N2454_0 ( .fault(fault), .net(N2454), .FEN(FEN[1167]), .op(N2454_t0) );
fim FAN_N2454_1 ( .fault(fault), .net(N2454), .FEN(FEN[1168]), .op(N2454_t1) );
fim FAN_N2454_2 ( .fault(fault), .net(N2454), .FEN(FEN[1169]), .op(N2454_t2) );
fim FAN_N2662_0 ( .fault(fault), .net(N2662), .FEN(FEN[1170]), .op(N2662_t0) );
fim FAN_N2662_1 ( .fault(fault), .net(N2662), .FEN(FEN[1171]), .op(N2662_t1) );
fim FAN_N2662_2 ( .fault(fault), .net(N2662), .FEN(FEN[1172]), .op(N2662_t2) );
fim FAN_N2450_0 ( .fault(fault), .net(N2450), .FEN(FEN[1173]), .op(N2450_t0) );
fim FAN_N2450_1 ( .fault(fault), .net(N2450), .FEN(FEN[1174]), .op(N2450_t1) );
fim FAN_N2450_2 ( .fault(fault), .net(N2450), .FEN(FEN[1175]), .op(N2450_t2) );
fim FAN_N2658_0 ( .fault(fault), .net(N2658), .FEN(FEN[1176]), .op(N2658_t0) );
fim FAN_N2658_1 ( .fault(fault), .net(N2658), .FEN(FEN[1177]), .op(N2658_t1) );
fim FAN_N2658_2 ( .fault(fault), .net(N2658), .FEN(FEN[1178]), .op(N2658_t2) );
fim FAN_N2446_0 ( .fault(fault), .net(N2446), .FEN(FEN[1179]), .op(N2446_t0) );
fim FAN_N2446_1 ( .fault(fault), .net(N2446), .FEN(FEN[1180]), .op(N2446_t1) );
fim FAN_N2446_2 ( .fault(fault), .net(N2446), .FEN(FEN[1181]), .op(N2446_t2) );
fim FAN_N2654_0 ( .fault(fault), .net(N2654), .FEN(FEN[1182]), .op(N2654_t0) );
fim FAN_N2654_1 ( .fault(fault), .net(N2654), .FEN(FEN[1183]), .op(N2654_t1) );
fim FAN_N2654_2 ( .fault(fault), .net(N2654), .FEN(FEN[1184]), .op(N2654_t2) );
fim FAN_N2442_0 ( .fault(fault), .net(N2442), .FEN(FEN[1185]), .op(N2442_t0) );
fim FAN_N2442_1 ( .fault(fault), .net(N2442), .FEN(FEN[1186]), .op(N2442_t1) );
fim FAN_N2442_2 ( .fault(fault), .net(N2442), .FEN(FEN[1187]), .op(N2442_t2) );
fim FAN_N2650_0 ( .fault(fault), .net(N2650), .FEN(FEN[1188]), .op(N2650_t0) );
fim FAN_N2650_1 ( .fault(fault), .net(N2650), .FEN(FEN[1189]), .op(N2650_t1) );
fim FAN_N2781_0 ( .fault(fault), .net(N2781), .FEN(FEN[1190]), .op(N2781_t0) );
fim FAN_N2781_1 ( .fault(fault), .net(N2781), .FEN(FEN[1191]), .op(N2781_t1) );
fim FAN_N2604_0 ( .fault(fault), .net(N2604), .FEN(FEN[1192]), .op(N2604_t0) );
fim FAN_N2604_1 ( .fault(fault), .net(N2604), .FEN(FEN[1193]), .op(N2604_t1) );
fim FAN_N2790_0 ( .fault(fault), .net(N2790), .FEN(FEN[1194]), .op(N2790_t0) );
fim FAN_N2790_1 ( .fault(fault), .net(N2790), .FEN(FEN[1195]), .op(N2790_t1) );
fim FAN_N2793_0 ( .fault(fault), .net(N2793), .FEN(FEN[1196]), .op(N2793_t0) );
fim FAN_N2793_1 ( .fault(fault), .net(N2793), .FEN(FEN[1197]), .op(N2793_t1) );
fim FAN_N2796_0 ( .fault(fault), .net(N2796), .FEN(FEN[1198]), .op(N2796_t0) );
fim FAN_N2796_1 ( .fault(fault), .net(N2796), .FEN(FEN[1199]), .op(N2796_t1) );
fim FAN_N2766_0 ( .fault(fault), .net(N2766), .FEN(FEN[1200]), .op(N2766_t0) );
fim FAN_N2766_1 ( .fault(fault), .net(N2766), .FEN(FEN[1201]), .op(N2766_t1) );
fim FAN_N2769_0 ( .fault(fault), .net(N2769), .FEN(FEN[1202]), .op(N2769_t0) );
fim FAN_N2769_1 ( .fault(fault), .net(N2769), .FEN(FEN[1203]), .op(N2769_t1) );
fim FAN_N2772_0 ( .fault(fault), .net(N2772), .FEN(FEN[1204]), .op(N2772_t0) );
fim FAN_N2772_1 ( .fault(fault), .net(N2772), .FEN(FEN[1205]), .op(N2772_t1) );
fim FAN_N2775_0 ( .fault(fault), .net(N2775), .FEN(FEN[1206]), .op(N2775_t0) );
fim FAN_N2775_1 ( .fault(fault), .net(N2775), .FEN(FEN[1207]), .op(N2775_t1) );
fim FAN_N2674_0 ( .fault(fault), .net(N2674), .FEN(FEN[1208]), .op(N2674_t0) );
fim FAN_N2674_1 ( .fault(fault), .net(N2674), .FEN(FEN[1209]), .op(N2674_t1) );
fim FAN_N2674_2 ( .fault(fault), .net(N2674), .FEN(FEN[1210]), .op(N2674_t2) );
fim FAN_N2674_3 ( .fault(fault), .net(N2674), .FEN(FEN[1211]), .op(N2674_t3) );
fim FAN_N2674_4 ( .fault(fault), .net(N2674), .FEN(FEN[1212]), .op(N2674_t4) );
fim FAN_N2704_0 ( .fault(fault), .net(N2704), .FEN(FEN[1213]), .op(N2704_t0) );
fim FAN_N2704_1 ( .fault(fault), .net(N2704), .FEN(FEN[1214]), .op(N2704_t1) );
fim FAN_N2704_2 ( .fault(fault), .net(N2704), .FEN(FEN[1215]), .op(N2704_t2) );
fim FAN_N2700_0 ( .fault(fault), .net(N2700), .FEN(FEN[1216]), .op(N2700_t0) );
fim FAN_N2700_1 ( .fault(fault), .net(N2700), .FEN(FEN[1217]), .op(N2700_t1) );
fim FAN_N2700_2 ( .fault(fault), .net(N2700), .FEN(FEN[1218]), .op(N2700_t2) );
fim FAN_N2696_0 ( .fault(fault), .net(N2696), .FEN(FEN[1219]), .op(N2696_t0) );
fim FAN_N2696_1 ( .fault(fault), .net(N2696), .FEN(FEN[1220]), .op(N2696_t1) );
fim FAN_N2696_2 ( .fault(fault), .net(N2696), .FEN(FEN[1221]), .op(N2696_t2) );
fim FAN_N2688_0 ( .fault(fault), .net(N2688), .FEN(FEN[1222]), .op(N2688_t0) );
fim FAN_N2688_1 ( .fault(fault), .net(N2688), .FEN(FEN[1223]), .op(N2688_t1) );
fim FAN_N2688_2 ( .fault(fault), .net(N2688), .FEN(FEN[1224]), .op(N2688_t2) );
fim FAN_N2692_0 ( .fault(fault), .net(N2692), .FEN(FEN[1225]), .op(N2692_t0) );
fim FAN_N2692_1 ( .fault(fault), .net(N2692), .FEN(FEN[1226]), .op(N2692_t1) );
fim FAN_N2692_2 ( .fault(fault), .net(N2692), .FEN(FEN[1227]), .op(N2692_t2) );
fim FAN_N2784_0 ( .fault(fault), .net(N2784), .FEN(FEN[1228]), .op(N2784_t0) );
fim FAN_N2784_1 ( .fault(fault), .net(N2784), .FEN(FEN[1229]), .op(N2784_t1) );
fim FAN_N2787_0 ( .fault(fault), .net(N2787), .FEN(FEN[1230]), .op(N2787_t0) );
fim FAN_N2787_1 ( .fault(fault), .net(N2787), .FEN(FEN[1231]), .op(N2787_t1) );
fim FAN_N2611_0 ( .fault(fault), .net(N2611), .FEN(FEN[1232]), .op(N2611_t0) );
fim FAN_N2611_1 ( .fault(fault), .net(N2611), .FEN(FEN[1233]), .op(N2611_t1) );
fim FAN_N2611_2 ( .fault(fault), .net(N2611), .FEN(FEN[1234]), .op(N2611_t2) );
fim FAN_N2607_0 ( .fault(fault), .net(N2607), .FEN(FEN[1235]), .op(N2607_t0) );
fim FAN_N2607_1 ( .fault(fault), .net(N2607), .FEN(FEN[1236]), .op(N2607_t1) );
fim FAN_N2607_2 ( .fault(fault), .net(N2607), .FEN(FEN[1237]), .op(N2607_t2) );
fim FAN_N2615_0 ( .fault(fault), .net(N2615), .FEN(FEN[1238]), .op(N2615_t0) );
fim FAN_N2615_1 ( .fault(fault), .net(N2615), .FEN(FEN[1239]), .op(N2615_t1) );
fim FAN_N2615_2 ( .fault(fault), .net(N2615), .FEN(FEN[1240]), .op(N2615_t2) );
fim FAN_N2680_0 ( .fault(fault), .net(N2680), .FEN(FEN[1241]), .op(N2680_t0) );
fim FAN_N2680_1 ( .fault(fault), .net(N2680), .FEN(FEN[1242]), .op(N2680_t1) );
fim FAN_N3067_0 ( .fault(fault), .net(N3067), .FEN(FEN[1243]), .op(N3067_t0) );
fim FAN_N3067_1 ( .fault(fault), .net(N3067), .FEN(FEN[1244]), .op(N3067_t1) );
fim FAN_N3070_0 ( .fault(fault), .net(N3070), .FEN(FEN[1245]), .op(N3070_t0) );
fim FAN_N3070_1 ( .fault(fault), .net(N3070), .FEN(FEN[1246]), .op(N3070_t1) );
fim FAN_N3073_0 ( .fault(fault), .net(N3073), .FEN(FEN[1247]), .op(N3073_t0) );
fim FAN_N3073_1 ( .fault(fault), .net(N3073), .FEN(FEN[1248]), .op(N3073_t1) );
fim FAN_N3080_0 ( .fault(fault), .net(N3080), .FEN(FEN[1249]), .op(N3080_t0) );
fim FAN_N3080_1 ( .fault(fault), .net(N3080), .FEN(FEN[1250]), .op(N3080_t1) );
fim FAN_N3061_0 ( .fault(fault), .net(N3061), .FEN(FEN[1251]), .op(N3061_t0) );
fim FAN_N3061_1 ( .fault(fault), .net(N3061), .FEN(FEN[1252]), .op(N3061_t1) );
fim FAN_N3064_0 ( .fault(fault), .net(N3064), .FEN(FEN[1253]), .op(N3064_t0) );
fim FAN_N3064_1 ( .fault(fault), .net(N3064), .FEN(FEN[1254]), .op(N3064_t1) );
fim FAN_N3487_0 ( .fault(fault), .net(N3487), .FEN(FEN[1255]), .op(N3487_t0) );
fim FAN_N3487_1 ( .fault(fault), .net(N3487), .FEN(FEN[1256]), .op(N3487_t1) );
fim FAN_N3490_0 ( .fault(fault), .net(N3490), .FEN(FEN[1257]), .op(N3490_t0) );
fim FAN_N3490_1 ( .fault(fault), .net(N3490), .FEN(FEN[1258]), .op(N3490_t1) );
fim FAN_N3493_0 ( .fault(fault), .net(N3493), .FEN(FEN[1259]), .op(N3493_t0) );
fim FAN_N3493_1 ( .fault(fault), .net(N3493), .FEN(FEN[1260]), .op(N3493_t1) );
fim FAN_N3496_0 ( .fault(fault), .net(N3496), .FEN(FEN[1261]), .op(N3496_t0) );
fim FAN_N3496_1 ( .fault(fault), .net(N3496), .FEN(FEN[1262]), .op(N3496_t1) );
fim FAN_N3499_0 ( .fault(fault), .net(N3499), .FEN(FEN[1263]), .op(N3499_t0) );
fim FAN_N3499_1 ( .fault(fault), .net(N3499), .FEN(FEN[1264]), .op(N3499_t1) );
fim FAN_N3122_0 ( .fault(fault), .net(N3122), .FEN(FEN[1265]), .op(N3122_t0) );
fim FAN_N3122_1 ( .fault(fault), .net(N3122), .FEN(FEN[1266]), .op(N3122_t1) );
fim FAN_N3122_2 ( .fault(fault), .net(N3122), .FEN(FEN[1267]), .op(N3122_t2) );
fim FAN_N3126_0 ( .fault(fault), .net(N3126), .FEN(FEN[1268]), .op(N3126_t0) );
fim FAN_N3126_1 ( .fault(fault), .net(N3126), .FEN(FEN[1269]), .op(N3126_t1) );
fim FAN_N3126_2 ( .fault(fault), .net(N3126), .FEN(FEN[1270]), .op(N3126_t2) );
fim FAN_N3518_0 ( .fault(fault), .net(N3518), .FEN(FEN[1271]), .op(N3518_t0) );
fim FAN_N3518_1 ( .fault(fault), .net(N3518), .FEN(FEN[1272]), .op(N3518_t1) );
fim FAN_N3521_0 ( .fault(fault), .net(N3521), .FEN(FEN[1273]), .op(N3521_t0) );
fim FAN_N3521_1 ( .fault(fault), .net(N3521), .FEN(FEN[1274]), .op(N3521_t1) );
fim FAN_N3524_0 ( .fault(fault), .net(N3524), .FEN(FEN[1275]), .op(N3524_t0) );
fim FAN_N3524_1 ( .fault(fault), .net(N3524), .FEN(FEN[1276]), .op(N3524_t1) );
fim FAN_N3527_0 ( .fault(fault), .net(N3527), .FEN(FEN[1277]), .op(N3527_t0) );
fim FAN_N3527_1 ( .fault(fault), .net(N3527), .FEN(FEN[1278]), .op(N3527_t1) );
fim FAN_N3530_0 ( .fault(fault), .net(N3530), .FEN(FEN[1279]), .op(N3530_t0) );
fim FAN_N3530_1 ( .fault(fault), .net(N3530), .FEN(FEN[1280]), .op(N3530_t1) );
fim FAN_N3155_0 ( .fault(fault), .net(N3155), .FEN(FEN[1281]), .op(N3155_t0) );
fim FAN_N3155_1 ( .fault(fault), .net(N3155), .FEN(FEN[1282]), .op(N3155_t1) );
fim FAN_N3155_2 ( .fault(fault), .net(N3155), .FEN(FEN[1283]), .op(N3155_t2) );
fim FAN_N3159_0 ( .fault(fault), .net(N3159), .FEN(FEN[1284]), .op(N3159_t0) );
fim FAN_N3159_1 ( .fault(fault), .net(N3159), .FEN(FEN[1285]), .op(N3159_t1) );
fim FAN_N3159_2 ( .fault(fault), .net(N3159), .FEN(FEN[1286]), .op(N3159_t2) );
fim FAN_N3535_0 ( .fault(fault), .net(N3535), .FEN(FEN[1287]), .op(N3535_t0) );
fim FAN_N3535_1 ( .fault(fault), .net(N3535), .FEN(FEN[1288]), .op(N3535_t1) );
fim FAN_N3539_0 ( .fault(fault), .net(N3539), .FEN(FEN[1289]), .op(N3539_t0) );
fim FAN_N3539_1 ( .fault(fault), .net(N3539), .FEN(FEN[1290]), .op(N3539_t1) );
fim FAN_N3542_0 ( .fault(fault), .net(N3542), .FEN(FEN[1291]), .op(N3542_t0) );
fim FAN_N3542_1 ( .fault(fault), .net(N3542), .FEN(FEN[1292]), .op(N3542_t1) );
fim FAN_N3545_0 ( .fault(fault), .net(N3545), .FEN(FEN[1293]), .op(N3545_t0) );
fim FAN_N3545_1 ( .fault(fault), .net(N3545), .FEN(FEN[1294]), .op(N3545_t1) );
fim FAN_N3548_0 ( .fault(fault), .net(N3548), .FEN(FEN[1295]), .op(N3548_t0) );
fim FAN_N3548_1 ( .fault(fault), .net(N3548), .FEN(FEN[1296]), .op(N3548_t1) );
fim FAN_N3553_0 ( .fault(fault), .net(N3553), .FEN(FEN[1297]), .op(N3553_t0) );
fim FAN_N3553_1 ( .fault(fault), .net(N3553), .FEN(FEN[1298]), .op(N3553_t1) );
fim FAN_N3557_0 ( .fault(fault), .net(N3557), .FEN(FEN[1299]), .op(N3557_t0) );
fim FAN_N3557_1 ( .fault(fault), .net(N3557), .FEN(FEN[1300]), .op(N3557_t1) );
fim FAN_N3560_0 ( .fault(fault), .net(N3560), .FEN(FEN[1301]), .op(N3560_t0) );
fim FAN_N3560_1 ( .fault(fault), .net(N3560), .FEN(FEN[1302]), .op(N3560_t1) );
fim FAN_N3563_0 ( .fault(fault), .net(N3563), .FEN(FEN[1303]), .op(N3563_t0) );
fim FAN_N3563_1 ( .fault(fault), .net(N3563), .FEN(FEN[1304]), .op(N3563_t1) );
fim FAN_N3566_0 ( .fault(fault), .net(N3566), .FEN(FEN[1305]), .op(N3566_t0) );
fim FAN_N3566_1 ( .fault(fault), .net(N3566), .FEN(FEN[1306]), .op(N3566_t1) );
fim FAN_N3571_0 ( .fault(fault), .net(N3571), .FEN(FEN[1307]), .op(N3571_t0) );
fim FAN_N3571_1 ( .fault(fault), .net(N3571), .FEN(FEN[1308]), .op(N3571_t1) );
fim FAN_N3574_0 ( .fault(fault), .net(N3574), .FEN(FEN[1309]), .op(N3574_t0) );
fim FAN_N3574_1 ( .fault(fault), .net(N3574), .FEN(FEN[1310]), .op(N3574_t1) );
fim FAN_N3577_0 ( .fault(fault), .net(N3577), .FEN(FEN[1311]), .op(N3577_t0) );
fim FAN_N3577_1 ( .fault(fault), .net(N3577), .FEN(FEN[1312]), .op(N3577_t1) );
fim FAN_N3580_0 ( .fault(fault), .net(N3580), .FEN(FEN[1313]), .op(N3580_t0) );
fim FAN_N3580_1 ( .fault(fault), .net(N3580), .FEN(FEN[1314]), .op(N3580_t1) );
fim FAN_N3583_0 ( .fault(fault), .net(N3583), .FEN(FEN[1315]), .op(N3583_t0) );
fim FAN_N3583_1 ( .fault(fault), .net(N3583), .FEN(FEN[1316]), .op(N3583_t1) );
fim FAN_N3598_0 ( .fault(fault), .net(N3598), .FEN(FEN[1317]), .op(N3598_t0) );
fim FAN_N3598_1 ( .fault(fault), .net(N3598), .FEN(FEN[1318]), .op(N3598_t1) );
fim FAN_N3601_0 ( .fault(fault), .net(N3601), .FEN(FEN[1319]), .op(N3601_t0) );
fim FAN_N3601_1 ( .fault(fault), .net(N3601), .FEN(FEN[1320]), .op(N3601_t1) );
fim FAN_N3604_0 ( .fault(fault), .net(N3604), .FEN(FEN[1321]), .op(N3604_t0) );
fim FAN_N3604_1 ( .fault(fault), .net(N3604), .FEN(FEN[1322]), .op(N3604_t1) );
fim FAN_N3607_0 ( .fault(fault), .net(N3607), .FEN(FEN[1323]), .op(N3607_t0) );
fim FAN_N3607_1 ( .fault(fault), .net(N3607), .FEN(FEN[1324]), .op(N3607_t1) );
fim FAN_N3610_0 ( .fault(fault), .net(N3610), .FEN(FEN[1325]), .op(N3610_t0) );
fim FAN_N3610_1 ( .fault(fault), .net(N3610), .FEN(FEN[1326]), .op(N3610_t1) );
fim FAN_N3613_0 ( .fault(fault), .net(N3613), .FEN(FEN[1327]), .op(N3613_t0) );
fim FAN_N3613_1 ( .fault(fault), .net(N3613), .FEN(FEN[1328]), .op(N3613_t1) );
fim FAN_N3616_0 ( .fault(fault), .net(N3616), .FEN(FEN[1329]), .op(N3616_t0) );
fim FAN_N3616_1 ( .fault(fault), .net(N3616), .FEN(FEN[1330]), .op(N3616_t1) );
fim FAN_N3619_0 ( .fault(fault), .net(N3619), .FEN(FEN[1331]), .op(N3619_t0) );
fim FAN_N3619_1 ( .fault(fault), .net(N3619), .FEN(FEN[1332]), .op(N3619_t1) );
fim FAN_N3622_0 ( .fault(fault), .net(N3622), .FEN(FEN[1333]), .op(N3622_t0) );
fim FAN_N3622_1 ( .fault(fault), .net(N3622), .FEN(FEN[1334]), .op(N3622_t1) );
fim FAN_N3631_0 ( .fault(fault), .net(N3631), .FEN(FEN[1335]), .op(N3631_t0) );
fim FAN_N3631_1 ( .fault(fault), .net(N3631), .FEN(FEN[1336]), .op(N3631_t1) );
fim FAN_N3634_0 ( .fault(fault), .net(N3634), .FEN(FEN[1337]), .op(N3634_t0) );
fim FAN_N3634_1 ( .fault(fault), .net(N3634), .FEN(FEN[1338]), .op(N3634_t1) );
fim FAN_N3637_0 ( .fault(fault), .net(N3637), .FEN(FEN[1339]), .op(N3637_t0) );
fim FAN_N3637_1 ( .fault(fault), .net(N3637), .FEN(FEN[1340]), .op(N3637_t1) );
fim FAN_N3640_0 ( .fault(fault), .net(N3640), .FEN(FEN[1341]), .op(N3640_t0) );
fim FAN_N3640_1 ( .fault(fault), .net(N3640), .FEN(FEN[1342]), .op(N3640_t1) );
fim FAN_N3643_0 ( .fault(fault), .net(N3643), .FEN(FEN[1343]), .op(N3643_t0) );
fim FAN_N3643_1 ( .fault(fault), .net(N3643), .FEN(FEN[1344]), .op(N3643_t1) );
fim FAN_N3646_0 ( .fault(fault), .net(N3646), .FEN(FEN[1345]), .op(N3646_t0) );
fim FAN_N3646_1 ( .fault(fault), .net(N3646), .FEN(FEN[1346]), .op(N3646_t1) );
fim FAN_N3649_0 ( .fault(fault), .net(N3649), .FEN(FEN[1347]), .op(N3649_t0) );
fim FAN_N3649_1 ( .fault(fault), .net(N3649), .FEN(FEN[1348]), .op(N3649_t1) );
fim FAN_N3652_0 ( .fault(fault), .net(N3652), .FEN(FEN[1349]), .op(N3652_t0) );
fim FAN_N3652_1 ( .fault(fault), .net(N3652), .FEN(FEN[1350]), .op(N3652_t1) );
fim FAN_N3655_0 ( .fault(fault), .net(N3655), .FEN(FEN[1351]), .op(N3655_t0) );
fim FAN_N3655_1 ( .fault(fault), .net(N3655), .FEN(FEN[1352]), .op(N3655_t1) );
fim FAN_N3658_0 ( .fault(fault), .net(N3658), .FEN(FEN[1353]), .op(N3658_t0) );
fim FAN_N3658_1 ( .fault(fault), .net(N3658), .FEN(FEN[1354]), .op(N3658_t1) );
fim FAN_N3293_0 ( .fault(fault), .net(N3293), .FEN(FEN[1355]), .op(N3293_t0) );
fim FAN_N3293_1 ( .fault(fault), .net(N3293), .FEN(FEN[1356]), .op(N3293_t1) );
fim FAN_N3293_2 ( .fault(fault), .net(N3293), .FEN(FEN[1357]), .op(N3293_t2) );
fim FAN_N3293_3 ( .fault(fault), .net(N3293), .FEN(FEN[1358]), .op(N3293_t3) );
fim FAN_N3293_4 ( .fault(fault), .net(N3293), .FEN(FEN[1359]), .op(N3293_t4) );
fim FAN_N3287_0 ( .fault(fault), .net(N3287), .FEN(FEN[1360]), .op(N3287_t0) );
fim FAN_N3287_1 ( .fault(fault), .net(N3287), .FEN(FEN[1361]), .op(N3287_t1) );
fim FAN_N3287_2 ( .fault(fault), .net(N3287), .FEN(FEN[1362]), .op(N3287_t2) );
fim FAN_N3287_3 ( .fault(fault), .net(N3287), .FEN(FEN[1363]), .op(N3287_t3) );
fim FAN_N3287_4 ( .fault(fault), .net(N3287), .FEN(FEN[1364]), .op(N3287_t4) );
fim FAN_N3281_0 ( .fault(fault), .net(N3281), .FEN(FEN[1365]), .op(N3281_t0) );
fim FAN_N3281_1 ( .fault(fault), .net(N3281), .FEN(FEN[1366]), .op(N3281_t1) );
fim FAN_N3281_2 ( .fault(fault), .net(N3281), .FEN(FEN[1367]), .op(N3281_t2) );
fim FAN_N3281_3 ( .fault(fault), .net(N3281), .FEN(FEN[1368]), .op(N3281_t3) );
fim FAN_N3281_4 ( .fault(fault), .net(N3281), .FEN(FEN[1369]), .op(N3281_t4) );
fim FAN_N3273_0 ( .fault(fault), .net(N3273), .FEN(FEN[1370]), .op(N3273_t0) );
fim FAN_N3273_1 ( .fault(fault), .net(N3273), .FEN(FEN[1371]), .op(N3273_t1) );
fim FAN_N3273_2 ( .fault(fault), .net(N3273), .FEN(FEN[1372]), .op(N3273_t2) );
fim FAN_N3273_3 ( .fault(fault), .net(N3273), .FEN(FEN[1373]), .op(N3273_t3) );
fim FAN_N3273_4 ( .fault(fault), .net(N3273), .FEN(FEN[1374]), .op(N3273_t4) );
fim FAN_N3273_5 ( .fault(fault), .net(N3273), .FEN(FEN[1375]), .op(N3273_t5) );
fim FAN_N3273_6 ( .fault(fault), .net(N3273), .FEN(FEN[1376]), .op(N3273_t6) );
fim FAN_N3267_0 ( .fault(fault), .net(N3267), .FEN(FEN[1377]), .op(N3267_t0) );
fim FAN_N3267_1 ( .fault(fault), .net(N3267), .FEN(FEN[1378]), .op(N3267_t1) );
fim FAN_N3267_2 ( .fault(fault), .net(N3267), .FEN(FEN[1379]), .op(N3267_t2) );
fim FAN_N3267_3 ( .fault(fault), .net(N3267), .FEN(FEN[1380]), .op(N3267_t3) );
fim FAN_N3267_4 ( .fault(fault), .net(N3267), .FEN(FEN[1381]), .op(N3267_t4) );
fim FAN_N3355_0 ( .fault(fault), .net(N3355), .FEN(FEN[1382]), .op(N3355_t0) );
fim FAN_N3355_1 ( .fault(fault), .net(N3355), .FEN(FEN[1383]), .op(N3355_t1) );
fim FAN_N3355_2 ( .fault(fault), .net(N3355), .FEN(FEN[1384]), .op(N3355_t2) );
fim FAN_N3355_3 ( .fault(fault), .net(N3355), .FEN(FEN[1385]), .op(N3355_t3) );
fim FAN_N3355_4 ( .fault(fault), .net(N3355), .FEN(FEN[1386]), .op(N3355_t4) );
fim FAN_N3349_0 ( .fault(fault), .net(N3349), .FEN(FEN[1387]), .op(N3349_t0) );
fim FAN_N3349_1 ( .fault(fault), .net(N3349), .FEN(FEN[1388]), .op(N3349_t1) );
fim FAN_N3349_2 ( .fault(fault), .net(N3349), .FEN(FEN[1389]), .op(N3349_t2) );
fim FAN_N3349_3 ( .fault(fault), .net(N3349), .FEN(FEN[1390]), .op(N3349_t3) );
fim FAN_N3349_4 ( .fault(fault), .net(N3349), .FEN(FEN[1391]), .op(N3349_t4) );
fim FAN_N3343_0 ( .fault(fault), .net(N3343), .FEN(FEN[1392]), .op(N3343_t0) );
fim FAN_N3343_1 ( .fault(fault), .net(N3343), .FEN(FEN[1393]), .op(N3343_t1) );
fim FAN_N3343_2 ( .fault(fault), .net(N3343), .FEN(FEN[1394]), .op(N3343_t2) );
fim FAN_N3343_3 ( .fault(fault), .net(N3343), .FEN(FEN[1395]), .op(N3343_t3) );
fim FAN_N3343_4 ( .fault(fault), .net(N3343), .FEN(FEN[1396]), .op(N3343_t4) );
fim FAN_N3661_0 ( .fault(fault), .net(N3661), .FEN(FEN[1397]), .op(N3661_t0) );
fim FAN_N3661_1 ( .fault(fault), .net(N3661), .FEN(FEN[1398]), .op(N3661_t1) );
fim FAN_N3664_0 ( .fault(fault), .net(N3664), .FEN(FEN[1399]), .op(N3664_t0) );
fim FAN_N3664_1 ( .fault(fault), .net(N3664), .FEN(FEN[1400]), .op(N3664_t1) );
fim FAN_N3667_0 ( .fault(fault), .net(N3667), .FEN(FEN[1401]), .op(N3667_t0) );
fim FAN_N3667_1 ( .fault(fault), .net(N3667), .FEN(FEN[1402]), .op(N3667_t1) );
fim FAN_N3670_0 ( .fault(fault), .net(N3670), .FEN(FEN[1403]), .op(N3670_t0) );
fim FAN_N3670_1 ( .fault(fault), .net(N3670), .FEN(FEN[1404]), .op(N3670_t1) );
fim FAN_N3673_0 ( .fault(fault), .net(N3673), .FEN(FEN[1405]), .op(N3673_t0) );
fim FAN_N3673_1 ( .fault(fault), .net(N3673), .FEN(FEN[1406]), .op(N3673_t1) );
fim FAN_N3676_0 ( .fault(fault), .net(N3676), .FEN(FEN[1407]), .op(N3676_t0) );
fim FAN_N3676_1 ( .fault(fault), .net(N3676), .FEN(FEN[1408]), .op(N3676_t1) );
fim FAN_N3679_0 ( .fault(fault), .net(N3679), .FEN(FEN[1409]), .op(N3679_t0) );
fim FAN_N3679_1 ( .fault(fault), .net(N3679), .FEN(FEN[1410]), .op(N3679_t1) );
fim FAN_N3682_0 ( .fault(fault), .net(N3682), .FEN(FEN[1411]), .op(N3682_t0) );
fim FAN_N3682_1 ( .fault(fault), .net(N3682), .FEN(FEN[1412]), .op(N3682_t1) );
fim FAN_N3685_0 ( .fault(fault), .net(N3685), .FEN(FEN[1413]), .op(N3685_t0) );
fim FAN_N3685_1 ( .fault(fault), .net(N3685), .FEN(FEN[1414]), .op(N3685_t1) );
fim FAN_N3688_0 ( .fault(fault), .net(N3688), .FEN(FEN[1415]), .op(N3688_t0) );
fim FAN_N3688_1 ( .fault(fault), .net(N3688), .FEN(FEN[1416]), .op(N3688_t1) );
fim FAN_N3691_0 ( .fault(fault), .net(N3691), .FEN(FEN[1417]), .op(N3691_t0) );
fim FAN_N3691_1 ( .fault(fault), .net(N3691), .FEN(FEN[1418]), .op(N3691_t1) );
fim FAN_N3694_0 ( .fault(fault), .net(N3694), .FEN(FEN[1419]), .op(N3694_t0) );
fim FAN_N3694_1 ( .fault(fault), .net(N3694), .FEN(FEN[1420]), .op(N3694_t1) );
fim FAN_N3697_0 ( .fault(fault), .net(N3697), .FEN(FEN[1421]), .op(N3697_t0) );
fim FAN_N3697_1 ( .fault(fault), .net(N3697), .FEN(FEN[1422]), .op(N3697_t1) );
fim FAN_N3700_0 ( .fault(fault), .net(N3700), .FEN(FEN[1423]), .op(N3700_t0) );
fim FAN_N3700_1 ( .fault(fault), .net(N3700), .FEN(FEN[1424]), .op(N3700_t1) );
fim FAN_N3703_0 ( .fault(fault), .net(N3703), .FEN(FEN[1425]), .op(N3703_t0) );
fim FAN_N3703_1 ( .fault(fault), .net(N3703), .FEN(FEN[1426]), .op(N3703_t1) );
fim FAN_N3706_0 ( .fault(fault), .net(N3706), .FEN(FEN[1427]), .op(N3706_t0) );
fim FAN_N3706_1 ( .fault(fault), .net(N3706), .FEN(FEN[1428]), .op(N3706_t1) );
fim FAN_N3709_0 ( .fault(fault), .net(N3709), .FEN(FEN[1429]), .op(N3709_t0) );
fim FAN_N3709_1 ( .fault(fault), .net(N3709), .FEN(FEN[1430]), .op(N3709_t1) );
fim FAN_N3712_0 ( .fault(fault), .net(N3712), .FEN(FEN[1431]), .op(N3712_t0) );
fim FAN_N3712_1 ( .fault(fault), .net(N3712), .FEN(FEN[1432]), .op(N3712_t1) );
fim FAN_N3715_0 ( .fault(fault), .net(N3715), .FEN(FEN[1433]), .op(N3715_t0) );
fim FAN_N3715_1 ( .fault(fault), .net(N3715), .FEN(FEN[1434]), .op(N3715_t1) );
fim FAN_N3718_0 ( .fault(fault), .net(N3718), .FEN(FEN[1435]), .op(N3718_t0) );
fim FAN_N3718_1 ( .fault(fault), .net(N3718), .FEN(FEN[1436]), .op(N3718_t1) );
fim FAN_N3721_0 ( .fault(fault), .net(N3721), .FEN(FEN[1437]), .op(N3721_t0) );
fim FAN_N3721_1 ( .fault(fault), .net(N3721), .FEN(FEN[1438]), .op(N3721_t1) );
fim FAN_N3448_0 ( .fault(fault), .net(N3448), .FEN(FEN[1439]), .op(N3448_t0) );
fim FAN_N3448_1 ( .fault(fault), .net(N3448), .FEN(FEN[1440]), .op(N3448_t1) );
fim FAN_N3448_2 ( .fault(fault), .net(N3448), .FEN(FEN[1441]), .op(N3448_t2) );
fim FAN_N3724_0 ( .fault(fault), .net(N3724), .FEN(FEN[1442]), .op(N3724_t0) );
fim FAN_N3724_1 ( .fault(fault), .net(N3724), .FEN(FEN[1443]), .op(N3724_t1) );
fim FAN_N3444_0 ( .fault(fault), .net(N3444), .FEN(FEN[1444]), .op(N3444_t0) );
fim FAN_N3444_1 ( .fault(fault), .net(N3444), .FEN(FEN[1445]), .op(N3444_t1) );
fim FAN_N3444_2 ( .fault(fault), .net(N3444), .FEN(FEN[1446]), .op(N3444_t2) );
fim FAN_N3727_0 ( .fault(fault), .net(N3727), .FEN(FEN[1447]), .op(N3727_t0) );
fim FAN_N3727_1 ( .fault(fault), .net(N3727), .FEN(FEN[1448]), .op(N3727_t1) );
fim FAN_N3440_0 ( .fault(fault), .net(N3440), .FEN(FEN[1449]), .op(N3440_t0) );
fim FAN_N3440_1 ( .fault(fault), .net(N3440), .FEN(FEN[1450]), .op(N3440_t1) );
fim FAN_N3440_2 ( .fault(fault), .net(N3440), .FEN(FEN[1451]), .op(N3440_t2) );
fim FAN_N3436_0 ( .fault(fault), .net(N3436), .FEN(FEN[1452]), .op(N3436_t0) );
fim FAN_N3436_1 ( .fault(fault), .net(N3436), .FEN(FEN[1453]), .op(N3436_t1) );
fim FAN_N3436_2 ( .fault(fault), .net(N3436), .FEN(FEN[1454]), .op(N3436_t2) );
fim FAN_N3730_0 ( .fault(fault), .net(N3730), .FEN(FEN[1455]), .op(N3730_t0) );
fim FAN_N3730_1 ( .fault(fault), .net(N3730), .FEN(FEN[1456]), .op(N3730_t1) );
fim FAN_N3432_0 ( .fault(fault), .net(N3432), .FEN(FEN[1457]), .op(N3432_t0) );
fim FAN_N3432_1 ( .fault(fault), .net(N3432), .FEN(FEN[1458]), .op(N3432_t1) );
fim FAN_N3432_2 ( .fault(fault), .net(N3432), .FEN(FEN[1459]), .op(N3432_t2) );
fim FAN_N3428_0 ( .fault(fault), .net(N3428), .FEN(FEN[1460]), .op(N3428_t0) );
fim FAN_N3428_1 ( .fault(fault), .net(N3428), .FEN(FEN[1461]), .op(N3428_t1) );
fim FAN_N3428_2 ( .fault(fault), .net(N3428), .FEN(FEN[1462]), .op(N3428_t2) );
fim FAN_N3311_0 ( .fault(fault), .net(N3311), .FEN(FEN[1463]), .op(N3311_t0) );
fim FAN_N3311_1 ( .fault(fault), .net(N3311), .FEN(FEN[1464]), .op(N3311_t1) );
fim FAN_N3311_2 ( .fault(fault), .net(N3311), .FEN(FEN[1465]), .op(N3311_t2) );
fim FAN_N3424_0 ( .fault(fault), .net(N3424), .FEN(FEN[1466]), .op(N3424_t0) );
fim FAN_N3424_1 ( .fault(fault), .net(N3424), .FEN(FEN[1467]), .op(N3424_t1) );
fim FAN_N3424_2 ( .fault(fault), .net(N3424), .FEN(FEN[1468]), .op(N3424_t2) );
fim FAN_N3307_0 ( .fault(fault), .net(N3307), .FEN(FEN[1469]), .op(N3307_t0) );
fim FAN_N3307_1 ( .fault(fault), .net(N3307), .FEN(FEN[1470]), .op(N3307_t1) );
fim FAN_N3307_2 ( .fault(fault), .net(N3307), .FEN(FEN[1471]), .op(N3307_t2) );
fim FAN_N3420_0 ( .fault(fault), .net(N3420), .FEN(FEN[1472]), .op(N3420_t0) );
fim FAN_N3420_1 ( .fault(fault), .net(N3420), .FEN(FEN[1473]), .op(N3420_t1) );
fim FAN_N3420_2 ( .fault(fault), .net(N3420), .FEN(FEN[1474]), .op(N3420_t2) );
fim FAN_N3303_0 ( .fault(fault), .net(N3303), .FEN(FEN[1475]), .op(N3303_t0) );
fim FAN_N3303_1 ( .fault(fault), .net(N3303), .FEN(FEN[1476]), .op(N3303_t1) );
fim FAN_N3303_2 ( .fault(fault), .net(N3303), .FEN(FEN[1477]), .op(N3303_t2) );
fim FAN_N3416_0 ( .fault(fault), .net(N3416), .FEN(FEN[1478]), .op(N3416_t0) );
fim FAN_N3416_1 ( .fault(fault), .net(N3416), .FEN(FEN[1479]), .op(N3416_t1) );
fim FAN_N3416_2 ( .fault(fault), .net(N3416), .FEN(FEN[1480]), .op(N3416_t2) );
fim FAN_N3299_0 ( .fault(fault), .net(N3299), .FEN(FEN[1481]), .op(N3299_t0) );
fim FAN_N3299_1 ( .fault(fault), .net(N3299), .FEN(FEN[1482]), .op(N3299_t1) );
fim FAN_N3299_2 ( .fault(fault), .net(N3299), .FEN(FEN[1483]), .op(N3299_t2) );
fim FAN_N3733_0 ( .fault(fault), .net(N3733), .FEN(FEN[1484]), .op(N3733_t0) );
fim FAN_N3733_1 ( .fault(fault), .net(N3733), .FEN(FEN[1485]), .op(N3733_t1) );
fim FAN_N3736_0 ( .fault(fault), .net(N3736), .FEN(FEN[1486]), .op(N3736_t0) );
fim FAN_N3736_1 ( .fault(fault), .net(N3736), .FEN(FEN[1487]), .op(N3736_t1) );
fim FAN_N3739_0 ( .fault(fault), .net(N3739), .FEN(FEN[1488]), .op(N3739_t0) );
fim FAN_N3739_1 ( .fault(fault), .net(N3739), .FEN(FEN[1489]), .op(N3739_t1) );
fim FAN_N3742_0 ( .fault(fault), .net(N3742), .FEN(FEN[1490]), .op(N3742_t0) );
fim FAN_N3742_1 ( .fault(fault), .net(N3742), .FEN(FEN[1491]), .op(N3742_t1) );
fim FAN_N3745_0 ( .fault(fault), .net(N3745), .FEN(FEN[1492]), .op(N3745_t0) );
fim FAN_N3745_1 ( .fault(fault), .net(N3745), .FEN(FEN[1493]), .op(N3745_t1) );
fim FAN_N3748_0 ( .fault(fault), .net(N3748), .FEN(FEN[1494]), .op(N3748_t0) );
fim FAN_N3748_1 ( .fault(fault), .net(N3748), .FEN(FEN[1495]), .op(N3748_t1) );
fim FAN_N3751_0 ( .fault(fault), .net(N3751), .FEN(FEN[1496]), .op(N3751_t0) );
fim FAN_N3751_1 ( .fault(fault), .net(N3751), .FEN(FEN[1497]), .op(N3751_t1) );
fim FAN_N3754_0 ( .fault(fault), .net(N3754), .FEN(FEN[1498]), .op(N3754_t0) );
fim FAN_N3754_1 ( .fault(fault), .net(N3754), .FEN(FEN[1499]), .op(N3754_t1) );
fim FAN_N3757_0 ( .fault(fault), .net(N3757), .FEN(FEN[1500]), .op(N3757_t0) );
fim FAN_N3757_1 ( .fault(fault), .net(N3757), .FEN(FEN[1501]), .op(N3757_t1) );
fim FAN_N3760_0 ( .fault(fault), .net(N3760), .FEN(FEN[1502]), .op(N3760_t0) );
fim FAN_N3760_1 ( .fault(fault), .net(N3760), .FEN(FEN[1503]), .op(N3760_t1) );
fim FAN_N3763_0 ( .fault(fault), .net(N3763), .FEN(FEN[1504]), .op(N3763_t0) );
fim FAN_N3763_1 ( .fault(fault), .net(N3763), .FEN(FEN[1505]), .op(N3763_t1) );
fim FAN_N3375_0 ( .fault(fault), .net(N3375), .FEN(FEN[1506]), .op(N3375_t0) );
fim FAN_N3375_1 ( .fault(fault), .net(N3375), .FEN(FEN[1507]), .op(N3375_t1) );
fim FAN_N3375_2 ( .fault(fault), .net(N3375), .FEN(FEN[1508]), .op(N3375_t2) );
fim FAN_N3410_0 ( .fault(fault), .net(N3410), .FEN(FEN[1509]), .op(N3410_t0) );
fim FAN_N3410_1 ( .fault(fault), .net(N3410), .FEN(FEN[1510]), .op(N3410_t1) );
fim FAN_N3410_2 ( .fault(fault), .net(N3410), .FEN(FEN[1511]), .op(N3410_t2) );
fim FAN_N3410_3 ( .fault(fault), .net(N3410), .FEN(FEN[1512]), .op(N3410_t3) );
fim FAN_N3410_4 ( .fault(fault), .net(N3410), .FEN(FEN[1513]), .op(N3410_t4) );
fim FAN_N3404_0 ( .fault(fault), .net(N3404), .FEN(FEN[1514]), .op(N3404_t0) );
fim FAN_N3404_1 ( .fault(fault), .net(N3404), .FEN(FEN[1515]), .op(N3404_t1) );
fim FAN_N3404_2 ( .fault(fault), .net(N3404), .FEN(FEN[1516]), .op(N3404_t2) );
fim FAN_N3404_3 ( .fault(fault), .net(N3404), .FEN(FEN[1517]), .op(N3404_t3) );
fim FAN_N3404_4 ( .fault(fault), .net(N3404), .FEN(FEN[1518]), .op(N3404_t4) );
fim FAN_N3398_0 ( .fault(fault), .net(N3398), .FEN(FEN[1519]), .op(N3398_t0) );
fim FAN_N3398_1 ( .fault(fault), .net(N3398), .FEN(FEN[1520]), .op(N3398_t1) );
fim FAN_N3398_2 ( .fault(fault), .net(N3398), .FEN(FEN[1521]), .op(N3398_t2) );
fim FAN_N3398_3 ( .fault(fault), .net(N3398), .FEN(FEN[1522]), .op(N3398_t3) );
fim FAN_N3398_4 ( .fault(fault), .net(N3398), .FEN(FEN[1523]), .op(N3398_t4) );
fim FAN_N3390_0 ( .fault(fault), .net(N3390), .FEN(FEN[1524]), .op(N3390_t0) );
fim FAN_N3390_1 ( .fault(fault), .net(N3390), .FEN(FEN[1525]), .op(N3390_t1) );
fim FAN_N3390_2 ( .fault(fault), .net(N3390), .FEN(FEN[1526]), .op(N3390_t2) );
fim FAN_N3390_3 ( .fault(fault), .net(N3390), .FEN(FEN[1527]), .op(N3390_t3) );
fim FAN_N3390_4 ( .fault(fault), .net(N3390), .FEN(FEN[1528]), .op(N3390_t4) );
fim FAN_N3390_5 ( .fault(fault), .net(N3390), .FEN(FEN[1529]), .op(N3390_t5) );
fim FAN_N3390_6 ( .fault(fault), .net(N3390), .FEN(FEN[1530]), .op(N3390_t6) );
fim FAN_N3384_0 ( .fault(fault), .net(N3384), .FEN(FEN[1531]), .op(N3384_t0) );
fim FAN_N3384_1 ( .fault(fault), .net(N3384), .FEN(FEN[1532]), .op(N3384_t1) );
fim FAN_N3384_2 ( .fault(fault), .net(N3384), .FEN(FEN[1533]), .op(N3384_t2) );
fim FAN_N3384_3 ( .fault(fault), .net(N3384), .FEN(FEN[1534]), .op(N3384_t3) );
fim FAN_N3384_4 ( .fault(fault), .net(N3384), .FEN(FEN[1535]), .op(N3384_t4) );
fim FAN_N3334_0 ( .fault(fault), .net(N3334), .FEN(FEN[1536]), .op(N3334_t0) );
fim FAN_N3334_1 ( .fault(fault), .net(N3334), .FEN(FEN[1537]), .op(N3334_t1) );
fim FAN_N3334_2 ( .fault(fault), .net(N3334), .FEN(FEN[1538]), .op(N3334_t2) );
fim FAN_N3334_3 ( .fault(fault), .net(N3334), .FEN(FEN[1539]), .op(N3334_t3) );
fim FAN_N3334_4 ( .fault(fault), .net(N3334), .FEN(FEN[1540]), .op(N3334_t4) );
fim FAN_N3328_0 ( .fault(fault), .net(N3328), .FEN(FEN[1541]), .op(N3328_t0) );
fim FAN_N3328_1 ( .fault(fault), .net(N3328), .FEN(FEN[1542]), .op(N3328_t1) );
fim FAN_N3328_2 ( .fault(fault), .net(N3328), .FEN(FEN[1543]), .op(N3328_t2) );
fim FAN_N3328_3 ( .fault(fault), .net(N3328), .FEN(FEN[1544]), .op(N3328_t3) );
fim FAN_N3328_4 ( .fault(fault), .net(N3328), .FEN(FEN[1545]), .op(N3328_t4) );
fim FAN_N3322_0 ( .fault(fault), .net(N3322), .FEN(FEN[1546]), .op(N3322_t0) );
fim FAN_N3322_1 ( .fault(fault), .net(N3322), .FEN(FEN[1547]), .op(N3322_t1) );
fim FAN_N3322_2 ( .fault(fault), .net(N3322), .FEN(FEN[1548]), .op(N3322_t2) );
fim FAN_N3322_3 ( .fault(fault), .net(N3322), .FEN(FEN[1549]), .op(N3322_t3) );
fim FAN_N3322_4 ( .fault(fault), .net(N3322), .FEN(FEN[1550]), .op(N3322_t4) );
fim FAN_N3315_0 ( .fault(fault), .net(N3315), .FEN(FEN[1551]), .op(N3315_t0) );
fim FAN_N3315_1 ( .fault(fault), .net(N3315), .FEN(FEN[1552]), .op(N3315_t1) );
fim FAN_N3315_2 ( .fault(fault), .net(N3315), .FEN(FEN[1553]), .op(N3315_t2) );
fim FAN_N3315_3 ( .fault(fault), .net(N3315), .FEN(FEN[1554]), .op(N3315_t3) );
fim FAN_N3315_4 ( .fault(fault), .net(N3315), .FEN(FEN[1555]), .op(N3315_t4) );
fim FAN_N3315_5 ( .fault(fault), .net(N3315), .FEN(FEN[1556]), .op(N3315_t5) );
fim FAN_N3766_0 ( .fault(fault), .net(N3766), .FEN(FEN[1557]), .op(N3766_t0) );
fim FAN_N3766_1 ( .fault(fault), .net(N3766), .FEN(FEN[1558]), .op(N3766_t1) );
fim FAN_N3769_0 ( .fault(fault), .net(N3769), .FEN(FEN[1559]), .op(N3769_t0) );
fim FAN_N3769_1 ( .fault(fault), .net(N3769), .FEN(FEN[1560]), .op(N3769_t1) );
fim FAN_N3772_0 ( .fault(fault), .net(N3772), .FEN(FEN[1561]), .op(N3772_t0) );
fim FAN_N3772_1 ( .fault(fault), .net(N3772), .FEN(FEN[1562]), .op(N3772_t1) );
fim FAN_N3775_0 ( .fault(fault), .net(N3775), .FEN(FEN[1563]), .op(N3775_t0) );
fim FAN_N3775_1 ( .fault(fault), .net(N3775), .FEN(FEN[1564]), .op(N3775_t1) );
fim FAN_N3778_0 ( .fault(fault), .net(N3778), .FEN(FEN[1565]), .op(N3778_t0) );
fim FAN_N3778_1 ( .fault(fault), .net(N3778), .FEN(FEN[1566]), .op(N3778_t1) );
fim FAN_N3783_0 ( .fault(fault), .net(N3783), .FEN(FEN[1567]), .op(N3783_t0) );
fim FAN_N3783_1 ( .fault(fault), .net(N3783), .FEN(FEN[1568]), .op(N3783_t1) );
fim FAN_N3786_0 ( .fault(fault), .net(N3786), .FEN(FEN[1569]), .op(N3786_t0) );
fim FAN_N3786_1 ( .fault(fault), .net(N3786), .FEN(FEN[1570]), .op(N3786_t1) );
fim FAN_N3789_0 ( .fault(fault), .net(N3789), .FEN(FEN[1571]), .op(N3789_t0) );
fim FAN_N3789_1 ( .fault(fault), .net(N3789), .FEN(FEN[1572]), .op(N3789_t1) );
fim FAN_N3792_0 ( .fault(fault), .net(N3792), .FEN(FEN[1573]), .op(N3792_t0) );
fim FAN_N3792_1 ( .fault(fault), .net(N3792), .FEN(FEN[1574]), .op(N3792_t1) );
fim FAN_N3807_0 ( .fault(fault), .net(N3807), .FEN(FEN[1575]), .op(N3807_t0) );
fim FAN_N3807_1 ( .fault(fault), .net(N3807), .FEN(FEN[1576]), .op(N3807_t1) );
fim FAN_N3810_0 ( .fault(fault), .net(N3810), .FEN(FEN[1577]), .op(N3810_t0) );
fim FAN_N3810_1 ( .fault(fault), .net(N3810), .FEN(FEN[1578]), .op(N3810_t1) );
fim FAN_N3813_0 ( .fault(fault), .net(N3813), .FEN(FEN[1579]), .op(N3813_t0) );
fim FAN_N3813_1 ( .fault(fault), .net(N3813), .FEN(FEN[1580]), .op(N3813_t1) );
fim FAN_N3816_0 ( .fault(fault), .net(N3816), .FEN(FEN[1581]), .op(N3816_t0) );
fim FAN_N3816_1 ( .fault(fault), .net(N3816), .FEN(FEN[1582]), .op(N3816_t1) );
fim FAN_N3819_0 ( .fault(fault), .net(N3819), .FEN(FEN[1583]), .op(N3819_t0) );
fim FAN_N3819_1 ( .fault(fault), .net(N3819), .FEN(FEN[1584]), .op(N3819_t1) );
fim FAN_N3822_0 ( .fault(fault), .net(N3822), .FEN(FEN[1585]), .op(N3822_t0) );
fim FAN_N3822_1 ( .fault(fault), .net(N3822), .FEN(FEN[1586]), .op(N3822_t1) );
fim FAN_N3825_0 ( .fault(fault), .net(N3825), .FEN(FEN[1587]), .op(N3825_t0) );
fim FAN_N3825_1 ( .fault(fault), .net(N3825), .FEN(FEN[1588]), .op(N3825_t1) );
fim FAN_N3828_0 ( .fault(fault), .net(N3828), .FEN(FEN[1589]), .op(N3828_t0) );
fim FAN_N3828_1 ( .fault(fault), .net(N3828), .FEN(FEN[1590]), .op(N3828_t1) );
fim FAN_N3831_0 ( .fault(fault), .net(N3831), .FEN(FEN[1591]), .op(N3831_t0) );
fim FAN_N3831_1 ( .fault(fault), .net(N3831), .FEN(FEN[1592]), .op(N3831_t1) );
fim FAN_N3482_0 ( .fault(fault), .net(N3482), .FEN(FEN[1593]), .op(N3482_t0) );
fim FAN_N3482_1 ( .fault(fault), .net(N3482), .FEN(FEN[1594]), .op(N3482_t1) );
fim FAN_N3482_2 ( .fault(fault), .net(N3482), .FEN(FEN[1595]), .op(N3482_t2) );
fim FAN_N3263_0 ( .fault(fault), .net(N3263), .FEN(FEN[1596]), .op(N3263_t0) );
fim FAN_N3263_1 ( .fault(fault), .net(N3263), .FEN(FEN[1597]), .op(N3263_t1) );
fim FAN_N3263_2 ( .fault(fault), .net(N3263), .FEN(FEN[1598]), .op(N3263_t2) );
fim FAN_N3478_0 ( .fault(fault), .net(N3478), .FEN(FEN[1599]), .op(N3478_t0) );
fim FAN_N3478_1 ( .fault(fault), .net(N3478), .FEN(FEN[1600]), .op(N3478_t1) );
fim FAN_N3478_2 ( .fault(fault), .net(N3478), .FEN(FEN[1601]), .op(N3478_t2) );
fim FAN_N3259_0 ( .fault(fault), .net(N3259), .FEN(FEN[1602]), .op(N3259_t0) );
fim FAN_N3259_1 ( .fault(fault), .net(N3259), .FEN(FEN[1603]), .op(N3259_t1) );
fim FAN_N3259_2 ( .fault(fault), .net(N3259), .FEN(FEN[1604]), .op(N3259_t2) );
fim FAN_N3474_0 ( .fault(fault), .net(N3474), .FEN(FEN[1605]), .op(N3474_t0) );
fim FAN_N3474_1 ( .fault(fault), .net(N3474), .FEN(FEN[1606]), .op(N3474_t1) );
fim FAN_N3474_2 ( .fault(fault), .net(N3474), .FEN(FEN[1607]), .op(N3474_t2) );
fim FAN_N3255_0 ( .fault(fault), .net(N3255), .FEN(FEN[1608]), .op(N3255_t0) );
fim FAN_N3255_1 ( .fault(fault), .net(N3255), .FEN(FEN[1609]), .op(N3255_t1) );
fim FAN_N3255_2 ( .fault(fault), .net(N3255), .FEN(FEN[1610]), .op(N3255_t2) );
fim FAN_N3470_0 ( .fault(fault), .net(N3470), .FEN(FEN[1611]), .op(N3470_t0) );
fim FAN_N3470_1 ( .fault(fault), .net(N3470), .FEN(FEN[1612]), .op(N3470_t1) );
fim FAN_N3470_2 ( .fault(fault), .net(N3470), .FEN(FEN[1613]), .op(N3470_t2) );
fim FAN_N3251_0 ( .fault(fault), .net(N3251), .FEN(FEN[1614]), .op(N3251_t0) );
fim FAN_N3251_1 ( .fault(fault), .net(N3251), .FEN(FEN[1615]), .op(N3251_t1) );
fim FAN_N3251_2 ( .fault(fault), .net(N3251), .FEN(FEN[1616]), .op(N3251_t2) );
fim FAN_N3466_0 ( .fault(fault), .net(N3466), .FEN(FEN[1617]), .op(N3466_t0) );
fim FAN_N3466_1 ( .fault(fault), .net(N3466), .FEN(FEN[1618]), .op(N3466_t1) );
fim FAN_N3466_2 ( .fault(fault), .net(N3466), .FEN(FEN[1619]), .op(N3466_t2) );
fim FAN_N3247_0 ( .fault(fault), .net(N3247), .FEN(FEN[1620]), .op(N3247_t0) );
fim FAN_N3247_1 ( .fault(fault), .net(N3247), .FEN(FEN[1621]), .op(N3247_t1) );
fim FAN_N3247_2 ( .fault(fault), .net(N3247), .FEN(FEN[1622]), .op(N3247_t2) );
fim FAN_N3846_0 ( .fault(fault), .net(N3846), .FEN(FEN[1623]), .op(N3846_t0) );
fim FAN_N3846_1 ( .fault(fault), .net(N3846), .FEN(FEN[1624]), .op(N3846_t1) );
fim FAN_N3462_0 ( .fault(fault), .net(N3462), .FEN(FEN[1625]), .op(N3462_t0) );
fim FAN_N3462_1 ( .fault(fault), .net(N3462), .FEN(FEN[1626]), .op(N3462_t1) );
fim FAN_N3462_2 ( .fault(fault), .net(N3462), .FEN(FEN[1627]), .op(N3462_t2) );
fim FAN_N3849_0 ( .fault(fault), .net(N3849), .FEN(FEN[1628]), .op(N3849_t0) );
fim FAN_N3849_1 ( .fault(fault), .net(N3849), .FEN(FEN[1629]), .op(N3849_t1) );
fim FAN_N3458_0 ( .fault(fault), .net(N3458), .FEN(FEN[1630]), .op(N3458_t0) );
fim FAN_N3458_1 ( .fault(fault), .net(N3458), .FEN(FEN[1631]), .op(N3458_t1) );
fim FAN_N3458_2 ( .fault(fault), .net(N3458), .FEN(FEN[1632]), .op(N3458_t2) );
fim FAN_N3852_0 ( .fault(fault), .net(N3852), .FEN(FEN[1633]), .op(N3852_t0) );
fim FAN_N3852_1 ( .fault(fault), .net(N3852), .FEN(FEN[1634]), .op(N3852_t1) );
fim FAN_N3454_0 ( .fault(fault), .net(N3454), .FEN(FEN[1635]), .op(N3454_t0) );
fim FAN_N3454_1 ( .fault(fault), .net(N3454), .FEN(FEN[1636]), .op(N3454_t1) );
fim FAN_N3454_2 ( .fault(fault), .net(N3454), .FEN(FEN[1637]), .op(N3454_t2) );
fim FAN_N3381_0 ( .fault(fault), .net(N3381), .FEN(FEN[1638]), .op(N3381_t0) );
fim FAN_N3381_1 ( .fault(fault), .net(N3381), .FEN(FEN[1639]), .op(N3381_t1) );
fim FAN_N3855_0 ( .fault(fault), .net(N3855), .FEN(FEN[1640]), .op(N3855_t0) );
fim FAN_N3855_1 ( .fault(fault), .net(N3855), .FEN(FEN[1641]), .op(N3855_t1) );
fim FAN_N3340_0 ( .fault(fault), .net(N3340), .FEN(FEN[1642]), .op(N3340_t0) );
fim FAN_N3340_1 ( .fault(fault), .net(N3340), .FEN(FEN[1643]), .op(N3340_t1) );
fim FAN_N3858_0 ( .fault(fault), .net(N3858), .FEN(FEN[1644]), .op(N3858_t0) );
fim FAN_N3858_1 ( .fault(fault), .net(N3858), .FEN(FEN[1645]), .op(N3858_t1) );
fim FAN_N3861_0 ( .fault(fault), .net(N3861), .FEN(FEN[1646]), .op(N3861_t0) );
fim FAN_N3861_1 ( .fault(fault), .net(N3861), .FEN(FEN[1647]), .op(N3861_t1) );
fim FAN_N3864_0 ( .fault(fault), .net(N3864), .FEN(FEN[1648]), .op(N3864_t0) );
fim FAN_N3864_1 ( .fault(fault), .net(N3864), .FEN(FEN[1649]), .op(N3864_t1) );
fim FAN_N3867_0 ( .fault(fault), .net(N3867), .FEN(FEN[1650]), .op(N3867_t0) );
fim FAN_N3867_1 ( .fault(fault), .net(N3867), .FEN(FEN[1651]), .op(N3867_t1) );
fim FAN_N3870_0 ( .fault(fault), .net(N3870), .FEN(FEN[1652]), .op(N3870_t0) );
fim FAN_N3870_1 ( .fault(fault), .net(N3870), .FEN(FEN[1653]), .op(N3870_t1) );
fim FAN_N3885_0 ( .fault(fault), .net(N3885), .FEN(FEN[1654]), .op(N3885_t0) );
fim FAN_N3885_1 ( .fault(fault), .net(N3885), .FEN(FEN[1655]), .op(N3885_t1) );
fim FAN_N3888_0 ( .fault(fault), .net(N3888), .FEN(FEN[1656]), .op(N3888_t0) );
fim FAN_N3888_1 ( .fault(fault), .net(N3888), .FEN(FEN[1657]), .op(N3888_t1) );
fim FAN_N3891_0 ( .fault(fault), .net(N3891), .FEN(FEN[1658]), .op(N3891_t0) );
fim FAN_N3891_1 ( .fault(fault), .net(N3891), .FEN(FEN[1659]), .op(N3891_t1) );
fim FAN_N3131_0 ( .fault(fault), .net(N3131), .FEN(FEN[1660]), .op(N3131_t0) );
fim FAN_N3131_1 ( .fault(fault), .net(N3131), .FEN(FEN[1661]), .op(N3131_t1) );
fim FAN_N3502_0 ( .fault(fault), .net(N3502), .FEN(FEN[1662]), .op(N3502_t0) );
fim FAN_N3502_1 ( .fault(fault), .net(N3502), .FEN(FEN[1663]), .op(N3502_t1) );
fim FAN_N3507_0 ( .fault(fault), .net(N3507), .FEN(FEN[1664]), .op(N3507_t0) );
fim FAN_N3507_1 ( .fault(fault), .net(N3507), .FEN(FEN[1665]), .op(N3507_t1) );
fim FAN_N3510_0 ( .fault(fault), .net(N3510), .FEN(FEN[1666]), .op(N3510_t0) );
fim FAN_N3510_1 ( .fault(fault), .net(N3510), .FEN(FEN[1667]), .op(N3510_t1) );
fim FAN_N3515_0 ( .fault(fault), .net(N3515), .FEN(FEN[1668]), .op(N3515_t0) );
fim FAN_N3515_1 ( .fault(fault), .net(N3515), .FEN(FEN[1669]), .op(N3515_t1) );
fim FAN_N3114_0 ( .fault(fault), .net(N3114), .FEN(FEN[1670]), .op(N3114_t0) );
fim FAN_N3114_1 ( .fault(fault), .net(N3114), .FEN(FEN[1671]), .op(N3114_t1) );
fim FAN_N3114_2 ( .fault(fault), .net(N3114), .FEN(FEN[1672]), .op(N3114_t2) );
fim FAN_N3114_3 ( .fault(fault), .net(N3114), .FEN(FEN[1673]), .op(N3114_t3) );
fim FAN_N3114_4 ( .fault(fault), .net(N3114), .FEN(FEN[1674]), .op(N3114_t4) );
fim FAN_N3114_5 ( .fault(fault), .net(N3114), .FEN(FEN[1675]), .op(N3114_t5) );
fim FAN_N3114_6 ( .fault(fault), .net(N3114), .FEN(FEN[1676]), .op(N3114_t6) );
fim FAN_N3586_0 ( .fault(fault), .net(N3586), .FEN(FEN[1677]), .op(N3586_t0) );
fim FAN_N3586_1 ( .fault(fault), .net(N3586), .FEN(FEN[1678]), .op(N3586_t1) );
fim FAN_N3589_0 ( .fault(fault), .net(N3589), .FEN(FEN[1679]), .op(N3589_t0) );
fim FAN_N3589_1 ( .fault(fault), .net(N3589), .FEN(FEN[1680]), .op(N3589_t1) );
fim FAN_N3592_0 ( .fault(fault), .net(N3592), .FEN(FEN[1681]), .op(N3592_t0) );
fim FAN_N3592_1 ( .fault(fault), .net(N3592), .FEN(FEN[1682]), .op(N3592_t1) );
fim FAN_N3595_0 ( .fault(fault), .net(N3595), .FEN(FEN[1683]), .op(N3595_t0) );
fim FAN_N3595_1 ( .fault(fault), .net(N3595), .FEN(FEN[1684]), .op(N3595_t1) );
fim FAN_N3625_0 ( .fault(fault), .net(N3625), .FEN(FEN[1685]), .op(N3625_t0) );
fim FAN_N3625_1 ( .fault(fault), .net(N3625), .FEN(FEN[1686]), .op(N3625_t1) );
fim FAN_N3178_0 ( .fault(fault), .net(N3178), .FEN(FEN[1687]), .op(N3178_t0) );
fim FAN_N3178_1 ( .fault(fault), .net(N3178), .FEN(FEN[1688]), .op(N3178_t1) );
fim FAN_N3178_2 ( .fault(fault), .net(N3178), .FEN(FEN[1689]), .op(N3178_t2) );
fim FAN_N3178_3 ( .fault(fault), .net(N3178), .FEN(FEN[1690]), .op(N3178_t3) );
fim FAN_N3178_4 ( .fault(fault), .net(N3178), .FEN(FEN[1691]), .op(N3178_t4) );
fim FAN_N3628_0 ( .fault(fault), .net(N3628), .FEN(FEN[1692]), .op(N3628_t0) );
fim FAN_N3628_1 ( .fault(fault), .net(N3628), .FEN(FEN[1693]), .op(N3628_t1) );
fim FAN_N3202_0 ( .fault(fault), .net(N3202), .FEN(FEN[1694]), .op(N3202_t0) );
fim FAN_N3202_1 ( .fault(fault), .net(N3202), .FEN(FEN[1695]), .op(N3202_t1) );
fim FAN_N3202_2 ( .fault(fault), .net(N3202), .FEN(FEN[1696]), .op(N3202_t2) );
fim FAN_N3202_3 ( .fault(fault), .net(N3202), .FEN(FEN[1697]), .op(N3202_t3) );
fim FAN_N3202_4 ( .fault(fault), .net(N3202), .FEN(FEN[1698]), .op(N3202_t4) );
fim FAN_N3202_5 ( .fault(fault), .net(N3202), .FEN(FEN[1699]), .op(N3202_t5) );
fim FAN_N3202_6 ( .fault(fault), .net(N3202), .FEN(FEN[1700]), .op(N3202_t6) );
fim FAN_N3221_0 ( .fault(fault), .net(N3221), .FEN(FEN[1701]), .op(N3221_t0) );
fim FAN_N3221_1 ( .fault(fault), .net(N3221), .FEN(FEN[1702]), .op(N3221_t1) );
fim FAN_N3221_2 ( .fault(fault), .net(N3221), .FEN(FEN[1703]), .op(N3221_t2) );
fim FAN_N3221_3 ( .fault(fault), .net(N3221), .FEN(FEN[1704]), .op(N3221_t3) );
fim FAN_N3221_4 ( .fault(fault), .net(N3221), .FEN(FEN[1705]), .op(N3221_t4) );
fim FAN_N3221_5 ( .fault(fault), .net(N3221), .FEN(FEN[1706]), .op(N3221_t5) );
fim FAN_N3795_0 ( .fault(fault), .net(N3795), .FEN(FEN[1707]), .op(N3795_t0) );
fim FAN_N3795_1 ( .fault(fault), .net(N3795), .FEN(FEN[1708]), .op(N3795_t1) );
fim FAN_N3798_0 ( .fault(fault), .net(N3798), .FEN(FEN[1709]), .op(N3798_t0) );
fim FAN_N3798_1 ( .fault(fault), .net(N3798), .FEN(FEN[1710]), .op(N3798_t1) );
fim FAN_N3801_0 ( .fault(fault), .net(N3801), .FEN(FEN[1711]), .op(N3801_t0) );
fim FAN_N3801_1 ( .fault(fault), .net(N3801), .FEN(FEN[1712]), .op(N3801_t1) );
fim FAN_N3804_0 ( .fault(fault), .net(N3804), .FEN(FEN[1713]), .op(N3804_t0) );
fim FAN_N3804_1 ( .fault(fault), .net(N3804), .FEN(FEN[1714]), .op(N3804_t1) );
fim FAN_N3834_0 ( .fault(fault), .net(N3834), .FEN(FEN[1715]), .op(N3834_t0) );
fim FAN_N3834_1 ( .fault(fault), .net(N3834), .FEN(FEN[1716]), .op(N3834_t1) );
fim FAN_N3837_0 ( .fault(fault), .net(N3837), .FEN(FEN[1717]), .op(N3837_t0) );
fim FAN_N3837_1 ( .fault(fault), .net(N3837), .FEN(FEN[1718]), .op(N3837_t1) );
fim FAN_N3840_0 ( .fault(fault), .net(N3840), .FEN(FEN[1719]), .op(N3840_t0) );
fim FAN_N3840_1 ( .fault(fault), .net(N3840), .FEN(FEN[1720]), .op(N3840_t1) );
fim FAN_N3843_0 ( .fault(fault), .net(N3843), .FEN(FEN[1721]), .op(N3843_t0) );
fim FAN_N3843_1 ( .fault(fault), .net(N3843), .FEN(FEN[1722]), .op(N3843_t1) );
fim FAN_N3873_0 ( .fault(fault), .net(N3873), .FEN(FEN[1723]), .op(N3873_t0) );
fim FAN_N3873_1 ( .fault(fault), .net(N3873), .FEN(FEN[1724]), .op(N3873_t1) );
fim FAN_N3876_0 ( .fault(fault), .net(N3876), .FEN(FEN[1725]), .op(N3876_t0) );
fim FAN_N3876_1 ( .fault(fault), .net(N3876), .FEN(FEN[1726]), .op(N3876_t1) );
fim FAN_N3879_0 ( .fault(fault), .net(N3879), .FEN(FEN[1727]), .op(N3879_t0) );
fim FAN_N3879_1 ( .fault(fault), .net(N3879), .FEN(FEN[1728]), .op(N3879_t1) );
fim FAN_N3882_0 ( .fault(fault), .net(N3882), .FEN(FEN[1729]), .op(N3882_t0) );
fim FAN_N3882_1 ( .fault(fault), .net(N3882), .FEN(FEN[1730]), .op(N3882_t1) );
fim FAN_N4193_0 ( .fault(fault), .net(N4193), .FEN(FEN[1731]), .op(N4193_t0) );
fim FAN_N4193_1 ( .fault(fault), .net(N4193), .FEN(FEN[1732]), .op(N4193_t1) );
fim FAN_N4193_2 ( .fault(fault), .net(N4193), .FEN(FEN[1733]), .op(N4193_t2) );
fim FAN_N4303_0 ( .fault(fault), .net(N4303), .FEN(FEN[1734]), .op(N4303_t0) );
fim FAN_N4303_1 ( .fault(fault), .net(N4303), .FEN(FEN[1735]), .op(N4303_t1) );
fim FAN_N4803_0 ( .fault(fault), .net(N4803), .FEN(FEN[1736]), .op(N4803_t0) );
fim FAN_N4803_1 ( .fault(fault), .net(N4803), .FEN(FEN[1737]), .op(N4803_t1) );
fim FAN_N4806_0 ( .fault(fault), .net(N4806), .FEN(FEN[1738]), .op(N4806_t0) );
fim FAN_N4806_1 ( .fault(fault), .net(N4806), .FEN(FEN[1739]), .op(N4806_t1) );
fim FAN_N4817_0 ( .fault(fault), .net(N4817), .FEN(FEN[1740]), .op(N4817_t0) );
fim FAN_N4817_1 ( .fault(fault), .net(N4817), .FEN(FEN[1741]), .op(N4817_t1) );
fim FAN_N4820_0 ( .fault(fault), .net(N4820), .FEN(FEN[1742]), .op(N4820_t0) );
fim FAN_N4820_1 ( .fault(fault), .net(N4820), .FEN(FEN[1743]), .op(N4820_t1) );
fim FAN_N4823_0 ( .fault(fault), .net(N4823), .FEN(FEN[1744]), .op(N4823_t0) );
fim FAN_N4823_1 ( .fault(fault), .net(N4823), .FEN(FEN[1745]), .op(N4823_t1) );
fim FAN_N4826_0 ( .fault(fault), .net(N4826), .FEN(FEN[1746]), .op(N4826_t0) );
fim FAN_N4826_1 ( .fault(fault), .net(N4826), .FEN(FEN[1747]), .op(N4826_t1) );
fim FAN_N4829_0 ( .fault(fault), .net(N4829), .FEN(FEN[1748]), .op(N4829_t0) );
fim FAN_N4829_1 ( .fault(fault), .net(N4829), .FEN(FEN[1749]), .op(N4829_t1) );
fim FAN_N4832_0 ( .fault(fault), .net(N4832), .FEN(FEN[1750]), .op(N4832_t0) );
fim FAN_N4832_1 ( .fault(fault), .net(N4832), .FEN(FEN[1751]), .op(N4832_t1) );
fim FAN_N4835_0 ( .fault(fault), .net(N4835), .FEN(FEN[1752]), .op(N4835_t0) );
fim FAN_N4835_1 ( .fault(fault), .net(N4835), .FEN(FEN[1753]), .op(N4835_t1) );
fim FAN_N4838_0 ( .fault(fault), .net(N4838), .FEN(FEN[1754]), .op(N4838_t0) );
fim FAN_N4838_1 ( .fault(fault), .net(N4838), .FEN(FEN[1755]), .op(N4838_t1) );
fim FAN_N4841_0 ( .fault(fault), .net(N4841), .FEN(FEN[1756]), .op(N4841_t0) );
fim FAN_N4841_1 ( .fault(fault), .net(N4841), .FEN(FEN[1757]), .op(N4841_t1) );
fim FAN_N4769_0 ( .fault(fault), .net(N4769), .FEN(FEN[1758]), .op(N4769_t0) );
fim FAN_N4769_1 ( .fault(fault), .net(N4769), .FEN(FEN[1759]), .op(N4769_t1) );
fim FAN_N4769_2 ( .fault(fault), .net(N4769), .FEN(FEN[1760]), .op(N4769_t2) );
fim FAN_N4769_3 ( .fault(fault), .net(N4769), .FEN(FEN[1761]), .op(N4769_t3) );
fim FAN_N4769_4 ( .fault(fault), .net(N4769), .FEN(FEN[1762]), .op(N4769_t4) );
fim FAN_N4844_0 ( .fault(fault), .net(N4844), .FEN(FEN[1763]), .op(N4844_t0) );
fim FAN_N4844_1 ( .fault(fault), .net(N4844), .FEN(FEN[1764]), .op(N4844_t1) );
fim FAN_N4847_0 ( .fault(fault), .net(N4847), .FEN(FEN[1765]), .op(N4847_t0) );
fim FAN_N4847_1 ( .fault(fault), .net(N4847), .FEN(FEN[1766]), .op(N4847_t1) );
fim FAN_N4850_0 ( .fault(fault), .net(N4850), .FEN(FEN[1767]), .op(N4850_t0) );
fim FAN_N4850_1 ( .fault(fault), .net(N4850), .FEN(FEN[1768]), .op(N4850_t1) );
fim FAN_N4853_0 ( .fault(fault), .net(N4853), .FEN(FEN[1769]), .op(N4853_t0) );
fim FAN_N4853_1 ( .fault(fault), .net(N4853), .FEN(FEN[1770]), .op(N4853_t1) );
fim FAN_N4856_0 ( .fault(fault), .net(N4856), .FEN(FEN[1771]), .op(N4856_t0) );
fim FAN_N4856_1 ( .fault(fault), .net(N4856), .FEN(FEN[1772]), .op(N4856_t1) );
fim FAN_N4859_0 ( .fault(fault), .net(N4859), .FEN(FEN[1773]), .op(N4859_t0) );
fim FAN_N4859_1 ( .fault(fault), .net(N4859), .FEN(FEN[1774]), .op(N4859_t1) );
fim FAN_N4862_0 ( .fault(fault), .net(N4862), .FEN(FEN[1775]), .op(N4862_t0) );
fim FAN_N4862_1 ( .fault(fault), .net(N4862), .FEN(FEN[1776]), .op(N4862_t1) );
fim FAN_N4865_0 ( .fault(fault), .net(N4865), .FEN(FEN[1777]), .op(N4865_t0) );
fim FAN_N4865_1 ( .fault(fault), .net(N4865), .FEN(FEN[1778]), .op(N4865_t1) );
fim FAN_N4868_0 ( .fault(fault), .net(N4868), .FEN(FEN[1779]), .op(N4868_t0) );
fim FAN_N4868_1 ( .fault(fault), .net(N4868), .FEN(FEN[1780]), .op(N4868_t1) );
fim FAN_N4874_0 ( .fault(fault), .net(N4874), .FEN(FEN[1781]), .op(N4874_t0) );
fim FAN_N4874_1 ( .fault(fault), .net(N4874), .FEN(FEN[1782]), .op(N4874_t1) );
fim FAN_N4877_0 ( .fault(fault), .net(N4877), .FEN(FEN[1783]), .op(N4877_t0) );
fim FAN_N4877_1 ( .fault(fault), .net(N4877), .FEN(FEN[1784]), .op(N4877_t1) );
fim FAN_N4880_0 ( .fault(fault), .net(N4880), .FEN(FEN[1785]), .op(N4880_t0) );
fim FAN_N4880_1 ( .fault(fault), .net(N4880), .FEN(FEN[1786]), .op(N4880_t1) );
fim FAN_N4883_0 ( .fault(fault), .net(N4883), .FEN(FEN[1787]), .op(N4883_t0) );
fim FAN_N4883_1 ( .fault(fault), .net(N4883), .FEN(FEN[1788]), .op(N4883_t1) );
fim FAN_N4886_0 ( .fault(fault), .net(N4886), .FEN(FEN[1789]), .op(N4886_t0) );
fim FAN_N4886_1 ( .fault(fault), .net(N4886), .FEN(FEN[1790]), .op(N4886_t1) );
fim FAN_N4889_0 ( .fault(fault), .net(N4889), .FEN(FEN[1791]), .op(N4889_t0) );
fim FAN_N4889_1 ( .fault(fault), .net(N4889), .FEN(FEN[1792]), .op(N4889_t1) );
fim FAN_N4892_0 ( .fault(fault), .net(N4892), .FEN(FEN[1793]), .op(N4892_t0) );
fim FAN_N4892_1 ( .fault(fault), .net(N4892), .FEN(FEN[1794]), .op(N4892_t1) );
fim FAN_N4895_0 ( .fault(fault), .net(N4895), .FEN(FEN[1795]), .op(N4895_t0) );
fim FAN_N4895_1 ( .fault(fault), .net(N4895), .FEN(FEN[1796]), .op(N4895_t1) );
fim FAN_N4898_0 ( .fault(fault), .net(N4898), .FEN(FEN[1797]), .op(N4898_t0) );
fim FAN_N4898_1 ( .fault(fault), .net(N4898), .FEN(FEN[1798]), .op(N4898_t1) );
fim FAN_N4901_0 ( .fault(fault), .net(N4901), .FEN(FEN[1799]), .op(N4901_t0) );
fim FAN_N4901_1 ( .fault(fault), .net(N4901), .FEN(FEN[1800]), .op(N4901_t1) );
fim FAN_N4904_0 ( .fault(fault), .net(N4904), .FEN(FEN[1801]), .op(N4904_t0) );
fim FAN_N4904_1 ( .fault(fault), .net(N4904), .FEN(FEN[1802]), .op(N4904_t1) );
fim FAN_N4907_0 ( .fault(fault), .net(N4907), .FEN(FEN[1803]), .op(N4907_t0) );
fim FAN_N4907_1 ( .fault(fault), .net(N4907), .FEN(FEN[1804]), .op(N4907_t1) );
fim FAN_N4910_0 ( .fault(fault), .net(N4910), .FEN(FEN[1805]), .op(N4910_t0) );
fim FAN_N4910_1 ( .fault(fault), .net(N4910), .FEN(FEN[1806]), .op(N4910_t1) );
fim FAN_N4913_0 ( .fault(fault), .net(N4913), .FEN(FEN[1807]), .op(N4913_t0) );
fim FAN_N4913_1 ( .fault(fault), .net(N4913), .FEN(FEN[1808]), .op(N4913_t1) );
fim FAN_N4916_0 ( .fault(fault), .net(N4916), .FEN(FEN[1809]), .op(N4916_t0) );
fim FAN_N4916_1 ( .fault(fault), .net(N4916), .FEN(FEN[1810]), .op(N4916_t1) );
fim FAN_N4919_0 ( .fault(fault), .net(N4919), .FEN(FEN[1811]), .op(N4919_t0) );
fim FAN_N4919_1 ( .fault(fault), .net(N4919), .FEN(FEN[1812]), .op(N4919_t1) );
fim FAN_N4922_0 ( .fault(fault), .net(N4922), .FEN(FEN[1813]), .op(N4922_t0) );
fim FAN_N4922_1 ( .fault(fault), .net(N4922), .FEN(FEN[1814]), .op(N4922_t1) );
fim FAN_N4925_0 ( .fault(fault), .net(N4925), .FEN(FEN[1815]), .op(N4925_t0) );
fim FAN_N4925_1 ( .fault(fault), .net(N4925), .FEN(FEN[1816]), .op(N4925_t1) );
fim FAN_N4928_0 ( .fault(fault), .net(N4928), .FEN(FEN[1817]), .op(N4928_t0) );
fim FAN_N4928_1 ( .fault(fault), .net(N4928), .FEN(FEN[1818]), .op(N4928_t1) );
fim FAN_N4931_0 ( .fault(fault), .net(N4931), .FEN(FEN[1819]), .op(N4931_t0) );
fim FAN_N4931_1 ( .fault(fault), .net(N4931), .FEN(FEN[1820]), .op(N4931_t1) );
fim FAN_N4934_0 ( .fault(fault), .net(N4934), .FEN(FEN[1821]), .op(N4934_t0) );
fim FAN_N4934_1 ( .fault(fault), .net(N4934), .FEN(FEN[1822]), .op(N4934_t1) );
fim FAN_N4937_0 ( .fault(fault), .net(N4937), .FEN(FEN[1823]), .op(N4937_t0) );
fim FAN_N4937_1 ( .fault(fault), .net(N4937), .FEN(FEN[1824]), .op(N4937_t1) );
fim FAN_N4940_0 ( .fault(fault), .net(N4940), .FEN(FEN[1825]), .op(N4940_t0) );
fim FAN_N4940_1 ( .fault(fault), .net(N4940), .FEN(FEN[1826]), .op(N4940_t1) );
fim FAN_N4943_0 ( .fault(fault), .net(N4943), .FEN(FEN[1827]), .op(N4943_t0) );
fim FAN_N4943_1 ( .fault(fault), .net(N4943), .FEN(FEN[1828]), .op(N4943_t1) );
fim FAN_N4946_0 ( .fault(fault), .net(N4946), .FEN(FEN[1829]), .op(N4946_t0) );
fim FAN_N4946_1 ( .fault(fault), .net(N4946), .FEN(FEN[1830]), .op(N4946_t1) );
fim FAN_N4949_0 ( .fault(fault), .net(N4949), .FEN(FEN[1831]), .op(N4949_t0) );
fim FAN_N4949_1 ( .fault(fault), .net(N4949), .FEN(FEN[1832]), .op(N4949_t1) );
fim FAN_N4952_0 ( .fault(fault), .net(N4952), .FEN(FEN[1833]), .op(N4952_t0) );
fim FAN_N4952_1 ( .fault(fault), .net(N4952), .FEN(FEN[1834]), .op(N4952_t1) );
fim FAN_N4955_0 ( .fault(fault), .net(N4955), .FEN(FEN[1835]), .op(N4955_t0) );
fim FAN_N4955_1 ( .fault(fault), .net(N4955), .FEN(FEN[1836]), .op(N4955_t1) );
fim FAN_N4970_0 ( .fault(fault), .net(N4970), .FEN(FEN[1837]), .op(N4970_t0) );
fim FAN_N4970_1 ( .fault(fault), .net(N4970), .FEN(FEN[1838]), .op(N4970_t1) );
fim FAN_N4973_0 ( .fault(fault), .net(N4973), .FEN(FEN[1839]), .op(N4973_t0) );
fim FAN_N4973_1 ( .fault(fault), .net(N4973), .FEN(FEN[1840]), .op(N4973_t1) );
fim FAN_N4976_0 ( .fault(fault), .net(N4976), .FEN(FEN[1841]), .op(N4976_t0) );
fim FAN_N4976_1 ( .fault(fault), .net(N4976), .FEN(FEN[1842]), .op(N4976_t1) );
fim FAN_N4979_0 ( .fault(fault), .net(N4979), .FEN(FEN[1843]), .op(N4979_t0) );
fim FAN_N4979_1 ( .fault(fault), .net(N4979), .FEN(FEN[1844]), .op(N4979_t1) );
fim FAN_N4982_0 ( .fault(fault), .net(N4982), .FEN(FEN[1845]), .op(N4982_t0) );
fim FAN_N4982_1 ( .fault(fault), .net(N4982), .FEN(FEN[1846]), .op(N4982_t1) );
fim FAN_N4997_0 ( .fault(fault), .net(N4997), .FEN(FEN[1847]), .op(N4997_t0) );
fim FAN_N4997_1 ( .fault(fault), .net(N4997), .FEN(FEN[1848]), .op(N4997_t1) );
fim FAN_N5000_0 ( .fault(fault), .net(N5000), .FEN(FEN[1849]), .op(N5000_t0) );
fim FAN_N5000_1 ( .fault(fault), .net(N5000), .FEN(FEN[1850]), .op(N5000_t1) );
fim FAN_N5003_0 ( .fault(fault), .net(N5003), .FEN(FEN[1851]), .op(N5003_t0) );
fim FAN_N5003_1 ( .fault(fault), .net(N5003), .FEN(FEN[1852]), .op(N5003_t1) );
fim FAN_N5006_0 ( .fault(fault), .net(N5006), .FEN(FEN[1853]), .op(N5006_t0) );
fim FAN_N5006_1 ( .fault(fault), .net(N5006), .FEN(FEN[1854]), .op(N5006_t1) );
fim FAN_N5009_0 ( .fault(fault), .net(N5009), .FEN(FEN[1855]), .op(N5009_t0) );
fim FAN_N5009_1 ( .fault(fault), .net(N5009), .FEN(FEN[1856]), .op(N5009_t1) );
fim FAN_N5012_0 ( .fault(fault), .net(N5012), .FEN(FEN[1857]), .op(N5012_t0) );
fim FAN_N5012_1 ( .fault(fault), .net(N5012), .FEN(FEN[1858]), .op(N5012_t1) );
fim FAN_N5015_0 ( .fault(fault), .net(N5015), .FEN(FEN[1859]), .op(N5015_t0) );
fim FAN_N5015_1 ( .fault(fault), .net(N5015), .FEN(FEN[1860]), .op(N5015_t1) );
fim FAN_N5018_0 ( .fault(fault), .net(N5018), .FEN(FEN[1861]), .op(N5018_t0) );
fim FAN_N5018_1 ( .fault(fault), .net(N5018), .FEN(FEN[1862]), .op(N5018_t1) );
fim FAN_N5021_0 ( .fault(fault), .net(N5021), .FEN(FEN[1863]), .op(N5021_t0) );
fim FAN_N5021_1 ( .fault(fault), .net(N5021), .FEN(FEN[1864]), .op(N5021_t1) );
fim FAN_N5024_0 ( .fault(fault), .net(N5024), .FEN(FEN[1865]), .op(N5024_t0) );
fim FAN_N5024_1 ( .fault(fault), .net(N5024), .FEN(FEN[1866]), .op(N5024_t1) );
fim FAN_N5033_0 ( .fault(fault), .net(N5033), .FEN(FEN[1867]), .op(N5033_t0) );
fim FAN_N5033_1 ( .fault(fault), .net(N5033), .FEN(FEN[1868]), .op(N5033_t1) );
fim FAN_N5036_0 ( .fault(fault), .net(N5036), .FEN(FEN[1869]), .op(N5036_t0) );
fim FAN_N5036_1 ( .fault(fault), .net(N5036), .FEN(FEN[1870]), .op(N5036_t1) );
fim FAN_N5039_0 ( .fault(fault), .net(N5039), .FEN(FEN[1871]), .op(N5039_t0) );
fim FAN_N5039_1 ( .fault(fault), .net(N5039), .FEN(FEN[1872]), .op(N5039_t1) );
fim FAN_N5042_0 ( .fault(fault), .net(N5042), .FEN(FEN[1873]), .op(N5042_t0) );
fim FAN_N5042_1 ( .fault(fault), .net(N5042), .FEN(FEN[1874]), .op(N5042_t1) );
fim FAN_N5049_0 ( .fault(fault), .net(N5049), .FEN(FEN[1875]), .op(N5049_t0) );
fim FAN_N5049_1 ( .fault(fault), .net(N5049), .FEN(FEN[1876]), .op(N5049_t1) );
fim FAN_N5068_0 ( .fault(fault), .net(N5068), .FEN(FEN[1877]), .op(N5068_t0) );
fim FAN_N5068_1 ( .fault(fault), .net(N5068), .FEN(FEN[1878]), .op(N5068_t1) );
fim FAN_N5071_0 ( .fault(fault), .net(N5071), .FEN(FEN[1879]), .op(N5071_t0) );
fim FAN_N5071_1 ( .fault(fault), .net(N5071), .FEN(FEN[1880]), .op(N5071_t1) );
fim FAN_N5074_0 ( .fault(fault), .net(N5074), .FEN(FEN[1881]), .op(N5074_t0) );
fim FAN_N5074_1 ( .fault(fault), .net(N5074), .FEN(FEN[1882]), .op(N5074_t1) );
fim FAN_N5077_0 ( .fault(fault), .net(N5077), .FEN(FEN[1883]), .op(N5077_t0) );
fim FAN_N5077_1 ( .fault(fault), .net(N5077), .FEN(FEN[1884]), .op(N5077_t1) );
fim FAN_N5080_0 ( .fault(fault), .net(N5080), .FEN(FEN[1885]), .op(N5080_t0) );
fim FAN_N5080_1 ( .fault(fault), .net(N5080), .FEN(FEN[1886]), .op(N5080_t1) );
fim FAN_N5083_0 ( .fault(fault), .net(N5083), .FEN(FEN[1887]), .op(N5083_t0) );
fim FAN_N5083_1 ( .fault(fault), .net(N5083), .FEN(FEN[1888]), .op(N5083_t1) );
fim FAN_N5086_0 ( .fault(fault), .net(N5086), .FEN(FEN[1889]), .op(N5086_t0) );
fim FAN_N5086_1 ( .fault(fault), .net(N5086), .FEN(FEN[1890]), .op(N5086_t1) );
fim FAN_N5089_0 ( .fault(fault), .net(N5089), .FEN(FEN[1891]), .op(N5089_t0) );
fim FAN_N5089_1 ( .fault(fault), .net(N5089), .FEN(FEN[1892]), .op(N5089_t1) );
fim FAN_N5092_0 ( .fault(fault), .net(N5092), .FEN(FEN[1893]), .op(N5092_t0) );
fim FAN_N5092_1 ( .fault(fault), .net(N5092), .FEN(FEN[1894]), .op(N5092_t1) );
fim FAN_N5095_0 ( .fault(fault), .net(N5095), .FEN(FEN[1895]), .op(N5095_t0) );
fim FAN_N5095_1 ( .fault(fault), .net(N5095), .FEN(FEN[1896]), .op(N5095_t1) );
fim FAN_N5098_0 ( .fault(fault), .net(N5098), .FEN(FEN[1897]), .op(N5098_t0) );
fim FAN_N5098_1 ( .fault(fault), .net(N5098), .FEN(FEN[1898]), .op(N5098_t1) );
fim FAN_N5101_0 ( .fault(fault), .net(N5101), .FEN(FEN[1899]), .op(N5101_t0) );
fim FAN_N5101_1 ( .fault(fault), .net(N5101), .FEN(FEN[1900]), .op(N5101_t1) );
fim FAN_N5104_0 ( .fault(fault), .net(N5104), .FEN(FEN[1901]), .op(N5104_t0) );
fim FAN_N5104_1 ( .fault(fault), .net(N5104), .FEN(FEN[1902]), .op(N5104_t1) );
fim FAN_N5107_0 ( .fault(fault), .net(N5107), .FEN(FEN[1903]), .op(N5107_t0) );
fim FAN_N5107_1 ( .fault(fault), .net(N5107), .FEN(FEN[1904]), .op(N5107_t1) );
fim FAN_N5114_0 ( .fault(fault), .net(N5114), .FEN(FEN[1905]), .op(N5114_t0) );
fim FAN_N5114_1 ( .fault(fault), .net(N5114), .FEN(FEN[1906]), .op(N5114_t1) );
fim FAN_N5117_0 ( .fault(fault), .net(N5117), .FEN(FEN[1907]), .op(N5117_t0) );
fim FAN_N5117_1 ( .fault(fault), .net(N5117), .FEN(FEN[1908]), .op(N5117_t1) );
fim FAN_N5120_0 ( .fault(fault), .net(N5120), .FEN(FEN[1909]), .op(N5120_t0) );
fim FAN_N5120_1 ( .fault(fault), .net(N5120), .FEN(FEN[1910]), .op(N5120_t1) );
fim FAN_N5123_0 ( .fault(fault), .net(N5123), .FEN(FEN[1911]), .op(N5123_t0) );
fim FAN_N5123_1 ( .fault(fault), .net(N5123), .FEN(FEN[1912]), .op(N5123_t1) );
fim FAN_N5138_0 ( .fault(fault), .net(N5138), .FEN(FEN[1913]), .op(N5138_t0) );
fim FAN_N5138_1 ( .fault(fault), .net(N5138), .FEN(FEN[1914]), .op(N5138_t1) );
fim FAN_N5141_0 ( .fault(fault), .net(N5141), .FEN(FEN[1915]), .op(N5141_t0) );
fim FAN_N5141_1 ( .fault(fault), .net(N5141), .FEN(FEN[1916]), .op(N5141_t1) );
fim FAN_N5144_0 ( .fault(fault), .net(N5144), .FEN(FEN[1917]), .op(N5144_t0) );
fim FAN_N5144_1 ( .fault(fault), .net(N5144), .FEN(FEN[1918]), .op(N5144_t1) );
fim FAN_N5147_0 ( .fault(fault), .net(N5147), .FEN(FEN[1919]), .op(N5147_t0) );
fim FAN_N5147_1 ( .fault(fault), .net(N5147), .FEN(FEN[1920]), .op(N5147_t1) );
fim FAN_N5150_0 ( .fault(fault), .net(N5150), .FEN(FEN[1921]), .op(N5150_t0) );
fim FAN_N5150_1 ( .fault(fault), .net(N5150), .FEN(FEN[1922]), .op(N5150_t1) );
fim FAN_N4784_0 ( .fault(fault), .net(N4784), .FEN(FEN[1923]), .op(N4784_t0) );
fim FAN_N4784_1 ( .fault(fault), .net(N4784), .FEN(FEN[1924]), .op(N4784_t1) );
fim FAN_N4790_0 ( .fault(fault), .net(N4790), .FEN(FEN[1925]), .op(N4790_t0) );
fim FAN_N4790_1 ( .fault(fault), .net(N4790), .FEN(FEN[1926]), .op(N4790_t1) );
fim FAN_N4796_0 ( .fault(fault), .net(N4796), .FEN(FEN[1927]), .op(N4796_t0) );
fim FAN_N4796_1 ( .fault(fault), .net(N4796), .FEN(FEN[1928]), .op(N4796_t1) );
fim FAN_N4810_0 ( .fault(fault), .net(N4810), .FEN(FEN[1929]), .op(N4810_t0) );
fim FAN_N4810_1 ( .fault(fault), .net(N4810), .FEN(FEN[1930]), .op(N4810_t1) );
fim FAN_N4814_0 ( .fault(fault), .net(N4814), .FEN(FEN[1931]), .op(N4814_t0) );
fim FAN_N4814_1 ( .fault(fault), .net(N4814), .FEN(FEN[1932]), .op(N4814_t1) );
fim FAN_N4555_0 ( .fault(fault), .net(N4555), .FEN(FEN[1933]), .op(N4555_t0) );
fim FAN_N4555_1 ( .fault(fault), .net(N4555), .FEN(FEN[1934]), .op(N4555_t1) );
fim FAN_N4555_2 ( .fault(fault), .net(N4555), .FEN(FEN[1935]), .op(N4555_t2) );
fim FAN_N4555_3 ( .fault(fault), .net(N4555), .FEN(FEN[1936]), .op(N4555_t3) );
fim FAN_N4555_4 ( .fault(fault), .net(N4555), .FEN(FEN[1937]), .op(N4555_t4) );
fim FAN_N4555_5 ( .fault(fault), .net(N4555), .FEN(FEN[1938]), .op(N4555_t5) );
fim FAN_N4871_0 ( .fault(fault), .net(N4871), .FEN(FEN[1939]), .op(N4871_t0) );
fim FAN_N4871_1 ( .fault(fault), .net(N4871), .FEN(FEN[1940]), .op(N4871_t1) );
fim FAN_N4586_0 ( .fault(fault), .net(N4586), .FEN(FEN[1941]), .op(N4586_t0) );
fim FAN_N4586_1 ( .fault(fault), .net(N4586), .FEN(FEN[1942]), .op(N4586_t1) );
fim FAN_N4586_2 ( .fault(fault), .net(N4586), .FEN(FEN[1943]), .op(N4586_t2) );
fim FAN_N4586_3 ( .fault(fault), .net(N4586), .FEN(FEN[1944]), .op(N4586_t3) );
fim FAN_N4586_4 ( .fault(fault), .net(N4586), .FEN(FEN[1945]), .op(N4586_t4) );
fim FAN_N4667_0 ( .fault(fault), .net(N4667), .FEN(FEN[1946]), .op(N4667_t0) );
fim FAN_N4667_1 ( .fault(fault), .net(N4667), .FEN(FEN[1947]), .op(N4667_t1) );
fim FAN_N4667_2 ( .fault(fault), .net(N4667), .FEN(FEN[1948]), .op(N4667_t2) );
fim FAN_N4667_3 ( .fault(fault), .net(N4667), .FEN(FEN[1949]), .op(N4667_t3) );
fim FAN_N4667_4 ( .fault(fault), .net(N4667), .FEN(FEN[1950]), .op(N4667_t4) );
fim FAN_N4667_5 ( .fault(fault), .net(N4667), .FEN(FEN[1951]), .op(N4667_t5) );
fim FAN_N4958_0 ( .fault(fault), .net(N4958), .FEN(FEN[1952]), .op(N4958_t0) );
fim FAN_N4958_1 ( .fault(fault), .net(N4958), .FEN(FEN[1953]), .op(N4958_t1) );
fim FAN_N4961_0 ( .fault(fault), .net(N4961), .FEN(FEN[1954]), .op(N4961_t0) );
fim FAN_N4961_1 ( .fault(fault), .net(N4961), .FEN(FEN[1955]), .op(N4961_t1) );
fim FAN_N4964_0 ( .fault(fault), .net(N4964), .FEN(FEN[1956]), .op(N4964_t0) );
fim FAN_N4964_1 ( .fault(fault), .net(N4964), .FEN(FEN[1957]), .op(N4964_t1) );
fim FAN_N4967_0 ( .fault(fault), .net(N4967), .FEN(FEN[1958]), .op(N4967_t0) );
fim FAN_N4967_1 ( .fault(fault), .net(N4967), .FEN(FEN[1959]), .op(N4967_t1) );
fim FAN_N4985_0 ( .fault(fault), .net(N4985), .FEN(FEN[1960]), .op(N4985_t0) );
fim FAN_N4985_1 ( .fault(fault), .net(N4985), .FEN(FEN[1961]), .op(N4985_t1) );
fim FAN_N4988_0 ( .fault(fault), .net(N4988), .FEN(FEN[1962]), .op(N4988_t0) );
fim FAN_N4988_1 ( .fault(fault), .net(N4988), .FEN(FEN[1963]), .op(N4988_t1) );
fim FAN_N4991_0 ( .fault(fault), .net(N4991), .FEN(FEN[1964]), .op(N4991_t0) );
fim FAN_N4991_1 ( .fault(fault), .net(N4991), .FEN(FEN[1965]), .op(N4991_t1) );
fim FAN_N4994_0 ( .fault(fault), .net(N4994), .FEN(FEN[1966]), .op(N4994_t0) );
fim FAN_N4994_1 ( .fault(fault), .net(N4994), .FEN(FEN[1967]), .op(N4994_t1) );
fim FAN_N5027_0 ( .fault(fault), .net(N5027), .FEN(FEN[1968]), .op(N5027_t0) );
fim FAN_N5027_1 ( .fault(fault), .net(N5027), .FEN(FEN[1969]), .op(N5027_t1) );
fim FAN_N4711_0 ( .fault(fault), .net(N4711), .FEN(FEN[1970]), .op(N4711_t0) );
fim FAN_N4711_1 ( .fault(fault), .net(N4711), .FEN(FEN[1971]), .op(N4711_t1) );
fim FAN_N4711_2 ( .fault(fault), .net(N4711), .FEN(FEN[1972]), .op(N4711_t2) );
fim FAN_N4711_3 ( .fault(fault), .net(N4711), .FEN(FEN[1973]), .op(N4711_t3) );
fim FAN_N4711_4 ( .fault(fault), .net(N4711), .FEN(FEN[1974]), .op(N4711_t4) );
fim FAN_N5030_0 ( .fault(fault), .net(N5030), .FEN(FEN[1975]), .op(N5030_t0) );
fim FAN_N5030_1 ( .fault(fault), .net(N5030), .FEN(FEN[1976]), .op(N5030_t1) );
fim FAN_N4735_0 ( .fault(fault), .net(N4735), .FEN(FEN[1977]), .op(N4735_t0) );
fim FAN_N4735_1 ( .fault(fault), .net(N4735), .FEN(FEN[1978]), .op(N4735_t1) );
fim FAN_N4735_2 ( .fault(fault), .net(N4735), .FEN(FEN[1979]), .op(N4735_t2) );
fim FAN_N4735_3 ( .fault(fault), .net(N4735), .FEN(FEN[1980]), .op(N4735_t3) );
fim FAN_N4735_4 ( .fault(fault), .net(N4735), .FEN(FEN[1981]), .op(N4735_t4) );
fim FAN_N4735_5 ( .fault(fault), .net(N4735), .FEN(FEN[1982]), .op(N4735_t5) );
fim FAN_N4735_6 ( .fault(fault), .net(N4735), .FEN(FEN[1983]), .op(N4735_t6) );
fim FAN_N5052_0 ( .fault(fault), .net(N5052), .FEN(FEN[1984]), .op(N5052_t0) );
fim FAN_N5052_1 ( .fault(fault), .net(N5052), .FEN(FEN[1985]), .op(N5052_t1) );
fim FAN_N5055_0 ( .fault(fault), .net(N5055), .FEN(FEN[1986]), .op(N5055_t0) );
fim FAN_N5055_1 ( .fault(fault), .net(N5055), .FEN(FEN[1987]), .op(N5055_t1) );
fim FAN_N5058_0 ( .fault(fault), .net(N5058), .FEN(FEN[1988]), .op(N5058_t0) );
fim FAN_N5058_1 ( .fault(fault), .net(N5058), .FEN(FEN[1989]), .op(N5058_t1) );
fim FAN_N5061_0 ( .fault(fault), .net(N5061), .FEN(FEN[1990]), .op(N5061_t0) );
fim FAN_N5061_1 ( .fault(fault), .net(N5061), .FEN(FEN[1991]), .op(N5061_t1) );
fim FAN_N5126_0 ( .fault(fault), .net(N5126), .FEN(FEN[1992]), .op(N5126_t0) );
fim FAN_N5126_1 ( .fault(fault), .net(N5126), .FEN(FEN[1993]), .op(N5126_t1) );
fim FAN_N5129_0 ( .fault(fault), .net(N5129), .FEN(FEN[1994]), .op(N5129_t0) );
fim FAN_N5129_1 ( .fault(fault), .net(N5129), .FEN(FEN[1995]), .op(N5129_t1) );
fim FAN_N5132_0 ( .fault(fault), .net(N5132), .FEN(FEN[1996]), .op(N5132_t0) );
fim FAN_N5132_1 ( .fault(fault), .net(N5132), .FEN(FEN[1997]), .op(N5132_t1) );
fim FAN_N5135_0 ( .fault(fault), .net(N5135), .FEN(FEN[1998]), .op(N5135_t0) );
fim FAN_N5135_1 ( .fault(fault), .net(N5135), .FEN(FEN[1999]), .op(N5135_t1) );
fim FAN_N5153_0 ( .fault(fault), .net(N5153), .FEN(FEN[2000]), .op(N5153_t0) );
fim FAN_N5153_1 ( .fault(fault), .net(N5153), .FEN(FEN[2001]), .op(N5153_t1) );
fim FAN_N5156_0 ( .fault(fault), .net(N5156), .FEN(FEN[2002]), .op(N5156_t0) );
fim FAN_N5156_1 ( .fault(fault), .net(N5156), .FEN(FEN[2003]), .op(N5156_t1) );
fim FAN_N5159_0 ( .fault(fault), .net(N5159), .FEN(FEN[2004]), .op(N5159_t0) );
fim FAN_N5159_1 ( .fault(fault), .net(N5159), .FEN(FEN[2005]), .op(N5159_t1) );
fim FAN_N5162_0 ( .fault(fault), .net(N5162), .FEN(FEN[2006]), .op(N5162_t0) );
fim FAN_N5162_1 ( .fault(fault), .net(N5162), .FEN(FEN[2007]), .op(N5162_t1) );
fim FAN_N5892_0 ( .fault(fault), .net(N5892), .FEN(FEN[2008]), .op(N5892_t0) );
fim FAN_N5892_1 ( .fault(fault), .net(N5892), .FEN(FEN[2009]), .op(N5892_t1) );
fim FAN_N5892_2 ( .fault(fault), .net(N5892), .FEN(FEN[2010]), .op(N5892_t2) );
fim FAN_N5892_3 ( .fault(fault), .net(N5892), .FEN(FEN[2011]), .op(N5892_t3) );
fim FAN_N5892_4 ( .fault(fault), .net(N5892), .FEN(FEN[2012]), .op(N5892_t4) );
fim FAN_N5683_0 ( .fault(fault), .net(N5683), .FEN(FEN[2013]), .op(N5683_t0) );
fim FAN_N5683_1 ( .fault(fault), .net(N5683), .FEN(FEN[2014]), .op(N5683_t1) );
fim FAN_N5683_2 ( .fault(fault), .net(N5683), .FEN(FEN[2015]), .op(N5683_t2) );
fim FAN_N5683_3 ( .fault(fault), .net(N5683), .FEN(FEN[2016]), .op(N5683_t3) );
fim FAN_N5683_4 ( .fault(fault), .net(N5683), .FEN(FEN[2017]), .op(N5683_t4) );
fim FAN_N5683_5 ( .fault(fault), .net(N5683), .FEN(FEN[2018]), .op(N5683_t5) );
fim FAN_N5670_0 ( .fault(fault), .net(N5670), .FEN(FEN[2019]), .op(N5670_t0) );
fim FAN_N5670_1 ( .fault(fault), .net(N5670), .FEN(FEN[2020]), .op(N5670_t1) );
fim FAN_N5670_2 ( .fault(fault), .net(N5670), .FEN(FEN[2021]), .op(N5670_t2) );
fim FAN_N5670_3 ( .fault(fault), .net(N5670), .FEN(FEN[2022]), .op(N5670_t3) );
fim FAN_N5670_4 ( .fault(fault), .net(N5670), .FEN(FEN[2023]), .op(N5670_t4) );
fim FAN_N5670_5 ( .fault(fault), .net(N5670), .FEN(FEN[2024]), .op(N5670_t5) );
fim FAN_N5670_6 ( .fault(fault), .net(N5670), .FEN(FEN[2025]), .op(N5670_t6) );
fim FAN_N5670_7 ( .fault(fault), .net(N5670), .FEN(FEN[2026]), .op(N5670_t7) );
fim FAN_N5670_8 ( .fault(fault), .net(N5670), .FEN(FEN[2027]), .op(N5670_t8) );
fim FAN_N5670_9 ( .fault(fault), .net(N5670), .FEN(FEN[2028]), .op(N5670_t9) );
fim FAN_N5670_10 ( .fault(fault), .net(N5670), .FEN(FEN[2029]), .op(N5670_t10) );
fim FAN_N5670_11 ( .fault(fault), .net(N5670), .FEN(FEN[2030]), .op(N5670_t11) );
fim FAN_N5654_0 ( .fault(fault), .net(N5654), .FEN(FEN[2031]), .op(N5654_t0) );
fim FAN_N5654_1 ( .fault(fault), .net(N5654), .FEN(FEN[2032]), .op(N5654_t1) );
fim FAN_N5654_2 ( .fault(fault), .net(N5654), .FEN(FEN[2033]), .op(N5654_t2) );
fim FAN_N5654_3 ( .fault(fault), .net(N5654), .FEN(FEN[2034]), .op(N5654_t3) );
fim FAN_N5654_4 ( .fault(fault), .net(N5654), .FEN(FEN[2035]), .op(N5654_t4) );
fim FAN_N5654_5 ( .fault(fault), .net(N5654), .FEN(FEN[2036]), .op(N5654_t5) );
fim FAN_N5654_6 ( .fault(fault), .net(N5654), .FEN(FEN[2037]), .op(N5654_t6) );
fim FAN_N5654_7 ( .fault(fault), .net(N5654), .FEN(FEN[2038]), .op(N5654_t7) );
fim FAN_N5654_8 ( .fault(fault), .net(N5654), .FEN(FEN[2039]), .op(N5654_t8) );
fim FAN_N5654_9 ( .fault(fault), .net(N5654), .FEN(FEN[2040]), .op(N5654_t9) );
fim FAN_N5654_10 ( .fault(fault), .net(N5654), .FEN(FEN[2041]), .op(N5654_t10) );
fim FAN_N5654_11 ( .fault(fault), .net(N5654), .FEN(FEN[2042]), .op(N5654_t11) );
fim FAN_N5654_12 ( .fault(fault), .net(N5654), .FEN(FEN[2043]), .op(N5654_t12) );
fim FAN_N5654_13 ( .fault(fault), .net(N5654), .FEN(FEN[2044]), .op(N5654_t13) );
fim FAN_N5654_14 ( .fault(fault), .net(N5654), .FEN(FEN[2045]), .op(N5654_t14) );
fim FAN_N5640_0 ( .fault(fault), .net(N5640), .FEN(FEN[2046]), .op(N5640_t0) );
fim FAN_N5640_1 ( .fault(fault), .net(N5640), .FEN(FEN[2047]), .op(N5640_t1) );
fim FAN_N5640_2 ( .fault(fault), .net(N5640), .FEN(FEN[2048]), .op(N5640_t2) );
fim FAN_N5640_3 ( .fault(fault), .net(N5640), .FEN(FEN[2049]), .op(N5640_t3) );
fim FAN_N5640_4 ( .fault(fault), .net(N5640), .FEN(FEN[2050]), .op(N5640_t4) );
fim FAN_N5640_5 ( .fault(fault), .net(N5640), .FEN(FEN[2051]), .op(N5640_t5) );
fim FAN_N5640_6 ( .fault(fault), .net(N5640), .FEN(FEN[2052]), .op(N5640_t6) );
fim FAN_N5640_7 ( .fault(fault), .net(N5640), .FEN(FEN[2053]), .op(N5640_t7) );
fim FAN_N5640_8 ( .fault(fault), .net(N5640), .FEN(FEN[2054]), .op(N5640_t8) );
fim FAN_N5640_9 ( .fault(fault), .net(N5640), .FEN(FEN[2055]), .op(N5640_t9) );
fim FAN_N5640_10 ( .fault(fault), .net(N5640), .FEN(FEN[2056]), .op(N5640_t10) );
fim FAN_N5640_11 ( .fault(fault), .net(N5640), .FEN(FEN[2057]), .op(N5640_t11) );
fim FAN_N5640_12 ( .fault(fault), .net(N5640), .FEN(FEN[2058]), .op(N5640_t12) );
fim FAN_N5632_0 ( .fault(fault), .net(N5632), .FEN(FEN[2059]), .op(N5632_t0) );
fim FAN_N5632_1 ( .fault(fault), .net(N5632), .FEN(FEN[2060]), .op(N5632_t1) );
fim FAN_N5632_2 ( .fault(fault), .net(N5632), .FEN(FEN[2061]), .op(N5632_t2) );
fim FAN_N5632_3 ( .fault(fault), .net(N5632), .FEN(FEN[2062]), .op(N5632_t3) );
fim FAN_N5632_4 ( .fault(fault), .net(N5632), .FEN(FEN[2063]), .op(N5632_t4) );
fim FAN_N5632_5 ( .fault(fault), .net(N5632), .FEN(FEN[2064]), .op(N5632_t5) );
fim FAN_N5632_6 ( .fault(fault), .net(N5632), .FEN(FEN[2065]), .op(N5632_t6) );
fim FAN_N3097_0 ( .fault(fault), .net(N3097), .FEN(FEN[2066]), .op(N3097_t0) );
fim FAN_N3097_1 ( .fault(fault), .net(N3097), .FEN(FEN[2067]), .op(N3097_t1) );
fim FAN_N3097_2 ( .fault(fault), .net(N3097), .FEN(FEN[2068]), .op(N3097_t2) );
fim FAN_N3101_0 ( .fault(fault), .net(N3101), .FEN(FEN[2069]), .op(N3101_t0) );
fim FAN_N3101_1 ( .fault(fault), .net(N3101), .FEN(FEN[2070]), .op(N3101_t1) );
fim FAN_N3101_2 ( .fault(fault), .net(N3101), .FEN(FEN[2071]), .op(N3101_t2) );
fim FAN_N3101_3 ( .fault(fault), .net(N3101), .FEN(FEN[2072]), .op(N3101_t3) );
fim FAN_N3101_4 ( .fault(fault), .net(N3101), .FEN(FEN[2073]), .op(N3101_t4) );
fim FAN_N3107_0 ( .fault(fault), .net(N3107), .FEN(FEN[2074]), .op(N3107_t0) );
fim FAN_N3107_1 ( .fault(fault), .net(N3107), .FEN(FEN[2075]), .op(N3107_t1) );
fim FAN_N3107_2 ( .fault(fault), .net(N3107), .FEN(FEN[2076]), .op(N3107_t2) );
fim FAN_N3107_3 ( .fault(fault), .net(N3107), .FEN(FEN[2077]), .op(N3107_t3) );
fim FAN_N3107_4 ( .fault(fault), .net(N3107), .FEN(FEN[2078]), .op(N3107_t4) );
fim FAN_N3107_5 ( .fault(fault), .net(N3107), .FEN(FEN[2079]), .op(N3107_t5) );
fim FAN_N5697_0 ( .fault(fault), .net(N5697), .FEN(FEN[2080]), .op(N5697_t0) );
fim FAN_N5697_1 ( .fault(fault), .net(N5697), .FEN(FEN[2081]), .op(N5697_t1) );
fim FAN_N5697_2 ( .fault(fault), .net(N5697), .FEN(FEN[2082]), .op(N5697_t2) );
fim FAN_N5697_3 ( .fault(fault), .net(N5697), .FEN(FEN[2083]), .op(N5697_t3) );
fim FAN_N5697_4 ( .fault(fault), .net(N5697), .FEN(FEN[2084]), .op(N5697_t4) );
fim FAN_N5697_5 ( .fault(fault), .net(N5697), .FEN(FEN[2085]), .op(N5697_t5) );
fim FAN_N5697_6 ( .fault(fault), .net(N5697), .FEN(FEN[2086]), .op(N5697_t6) );
fim FAN_N5697_7 ( .fault(fault), .net(N5697), .FEN(FEN[2087]), .op(N5697_t7) );
fim FAN_N5697_8 ( .fault(fault), .net(N5697), .FEN(FEN[2088]), .op(N5697_t8) );
fim FAN_N5728_0 ( .fault(fault), .net(N5728), .FEN(FEN[2089]), .op(N5728_t0) );
fim FAN_N5728_1 ( .fault(fault), .net(N5728), .FEN(FEN[2090]), .op(N5728_t1) );
fim FAN_N5728_2 ( .fault(fault), .net(N5728), .FEN(FEN[2091]), .op(N5728_t2) );
fim FAN_N5728_3 ( .fault(fault), .net(N5728), .FEN(FEN[2092]), .op(N5728_t3) );
fim FAN_N5728_4 ( .fault(fault), .net(N5728), .FEN(FEN[2093]), .op(N5728_t4) );
fim FAN_N5728_5 ( .fault(fault), .net(N5728), .FEN(FEN[2094]), .op(N5728_t5) );
fim FAN_N5707_0 ( .fault(fault), .net(N5707), .FEN(FEN[2095]), .op(N5707_t0) );
fim FAN_N5707_1 ( .fault(fault), .net(N5707), .FEN(FEN[2096]), .op(N5707_t1) );
fim FAN_N5707_2 ( .fault(fault), .net(N5707), .FEN(FEN[2097]), .op(N5707_t2) );
fim FAN_N5707_3 ( .fault(fault), .net(N5707), .FEN(FEN[2098]), .op(N5707_t3) );
fim FAN_N5707_4 ( .fault(fault), .net(N5707), .FEN(FEN[2099]), .op(N5707_t4) );
fim FAN_N5707_5 ( .fault(fault), .net(N5707), .FEN(FEN[2100]), .op(N5707_t5) );
fim FAN_N5707_6 ( .fault(fault), .net(N5707), .FEN(FEN[2101]), .op(N5707_t6) );
fim FAN_N5707_7 ( .fault(fault), .net(N5707), .FEN(FEN[2102]), .op(N5707_t7) );
fim FAN_N5707_8 ( .fault(fault), .net(N5707), .FEN(FEN[2103]), .op(N5707_t8) );
fim FAN_N5707_9 ( .fault(fault), .net(N5707), .FEN(FEN[2104]), .op(N5707_t9) );
fim FAN_N5690_0 ( .fault(fault), .net(N5690), .FEN(FEN[2105]), .op(N5690_t0) );
fim FAN_N5690_1 ( .fault(fault), .net(N5690), .FEN(FEN[2106]), .op(N5690_t1) );
fim FAN_N5690_2 ( .fault(fault), .net(N5690), .FEN(FEN[2107]), .op(N5690_t2) );
fim FAN_N5690_3 ( .fault(fault), .net(N5690), .FEN(FEN[2108]), .op(N5690_t3) );
fim FAN_N5690_4 ( .fault(fault), .net(N5690), .FEN(FEN[2109]), .op(N5690_t4) );
fim FAN_N5690_5 ( .fault(fault), .net(N5690), .FEN(FEN[2110]), .op(N5690_t5) );
fim FAN_N5718_0 ( .fault(fault), .net(N5718), .FEN(FEN[2111]), .op(N5718_t0) );
fim FAN_N5718_1 ( .fault(fault), .net(N5718), .FEN(FEN[2112]), .op(N5718_t1) );
fim FAN_N5718_2 ( .fault(fault), .net(N5718), .FEN(FEN[2113]), .op(N5718_t2) );
fim FAN_N5718_3 ( .fault(fault), .net(N5718), .FEN(FEN[2114]), .op(N5718_t3) );
fim FAN_N5718_4 ( .fault(fault), .net(N5718), .FEN(FEN[2115]), .op(N5718_t4) );
fim FAN_N5718_5 ( .fault(fault), .net(N5718), .FEN(FEN[2116]), .op(N5718_t5) );
fim FAN_N5718_6 ( .fault(fault), .net(N5718), .FEN(FEN[2117]), .op(N5718_t6) );
fim FAN_N5718_7 ( .fault(fault), .net(N5718), .FEN(FEN[2118]), .op(N5718_t7) );
fim FAN_N5718_8 ( .fault(fault), .net(N5718), .FEN(FEN[2119]), .op(N5718_t8) );
fim FAN_N3137_0 ( .fault(fault), .net(N3137), .FEN(FEN[2120]), .op(N3137_t0) );
fim FAN_N3137_1 ( .fault(fault), .net(N3137), .FEN(FEN[2121]), .op(N3137_t1) );
fim FAN_N3140_0 ( .fault(fault), .net(N3140), .FEN(FEN[2122]), .op(N3140_t0) );
fim FAN_N3140_1 ( .fault(fault), .net(N3140), .FEN(FEN[2123]), .op(N3140_t1) );
fim FAN_N3140_2 ( .fault(fault), .net(N3140), .FEN(FEN[2124]), .op(N3140_t2) );
fim FAN_N3144_0 ( .fault(fault), .net(N3144), .FEN(FEN[2125]), .op(N3144_t0) );
fim FAN_N3144_1 ( .fault(fault), .net(N3144), .FEN(FEN[2126]), .op(N3144_t1) );
fim FAN_N3144_2 ( .fault(fault), .net(N3144), .FEN(FEN[2127]), .op(N3144_t2) );
fim FAN_N3144_3 ( .fault(fault), .net(N3144), .FEN(FEN[2128]), .op(N3144_t3) );
fim FAN_N3149_0 ( .fault(fault), .net(N3149), .FEN(FEN[2129]), .op(N3149_t0) );
fim FAN_N3149_1 ( .fault(fault), .net(N3149), .FEN(FEN[2130]), .op(N3149_t1) );
fim FAN_N3149_2 ( .fault(fault), .net(N3149), .FEN(FEN[2131]), .op(N3149_t2) );
fim FAN_N3149_3 ( .fault(fault), .net(N3149), .FEN(FEN[2132]), .op(N3149_t3) );
fim FAN_N3149_4 ( .fault(fault), .net(N3149), .FEN(FEN[2133]), .op(N3149_t4) );
fim FAN_N5736_0 ( .fault(fault), .net(N5736), .FEN(FEN[2134]), .op(N5736_t0) );
fim FAN_N5736_1 ( .fault(fault), .net(N5736), .FEN(FEN[2135]), .op(N5736_t1) );
fim FAN_N5736_2 ( .fault(fault), .net(N5736), .FEN(FEN[2136]), .op(N5736_t2) );
fim FAN_N5740_0 ( .fault(fault), .net(N5740), .FEN(FEN[2137]), .op(N5740_t0) );
fim FAN_N5740_1 ( .fault(fault), .net(N5740), .FEN(FEN[2138]), .op(N5740_t1) );
fim FAN_N5740_2 ( .fault(fault), .net(N5740), .FEN(FEN[2139]), .op(N5740_t2) );
fim FAN_N5747_0 ( .fault(fault), .net(N5747), .FEN(FEN[2140]), .op(N5747_t0) );
fim FAN_N5747_1 ( .fault(fault), .net(N5747), .FEN(FEN[2141]), .op(N5747_t1) );
fim FAN_N5747_2 ( .fault(fault), .net(N5747), .FEN(FEN[2142]), .op(N5747_t2) );
fim FAN_N5751_0 ( .fault(fault), .net(N5751), .FEN(FEN[2143]), .op(N5751_t0) );
fim FAN_N5751_1 ( .fault(fault), .net(N5751), .FEN(FEN[2144]), .op(N5751_t1) );
fim FAN_N5751_2 ( .fault(fault), .net(N5751), .FEN(FEN[2145]), .op(N5751_t2) );
fim FAN_N5758_0 ( .fault(fault), .net(N5758), .FEN(FEN[2146]), .op(N5758_t0) );
fim FAN_N5758_1 ( .fault(fault), .net(N5758), .FEN(FEN[2147]), .op(N5758_t1) );
fim FAN_N5758_2 ( .fault(fault), .net(N5758), .FEN(FEN[2148]), .op(N5758_t2) );
fim FAN_N5762_0 ( .fault(fault), .net(N5762), .FEN(FEN[2149]), .op(N5762_t0) );
fim FAN_N5762_1 ( .fault(fault), .net(N5762), .FEN(FEN[2150]), .op(N5762_t1) );
fim FAN_N5762_2 ( .fault(fault), .net(N5762), .FEN(FEN[2151]), .op(N5762_t2) );
fim FAN_N5744_0 ( .fault(fault), .net(N5744), .FEN(FEN[2152]), .op(N5744_t0) );
fim FAN_N5744_1 ( .fault(fault), .net(N5744), .FEN(FEN[2153]), .op(N5744_t1) );
fim FAN_N5755_0 ( .fault(fault), .net(N5755), .FEN(FEN[2154]), .op(N5755_t0) );
fim FAN_N5755_1 ( .fault(fault), .net(N5755), .FEN(FEN[2155]), .op(N5755_t1) );
fim FAN_N5766_0 ( .fault(fault), .net(N5766), .FEN(FEN[2156]), .op(N5766_t0) );
fim FAN_N5766_1 ( .fault(fault), .net(N5766), .FEN(FEN[2157]), .op(N5766_t1) );
fim FAN_N5850_0 ( .fault(fault), .net(N5850), .FEN(FEN[2158]), .op(N5850_t0) );
fim FAN_N5850_1 ( .fault(fault), .net(N5850), .FEN(FEN[2159]), .op(N5850_t1) );
fim FAN_N5850_2 ( .fault(fault), .net(N5850), .FEN(FEN[2160]), .op(N5850_t2) );
fim FAN_N5850_3 ( .fault(fault), .net(N5850), .FEN(FEN[2161]), .op(N5850_t3) );
fim FAN_N5850_4 ( .fault(fault), .net(N5850), .FEN(FEN[2162]), .op(N5850_t4) );
fim FAN_N5789_0 ( .fault(fault), .net(N5789), .FEN(FEN[2163]), .op(N5789_t0) );
fim FAN_N5789_1 ( .fault(fault), .net(N5789), .FEN(FEN[2164]), .op(N5789_t1) );
fim FAN_N5789_2 ( .fault(fault), .net(N5789), .FEN(FEN[2165]), .op(N5789_t2) );
fim FAN_N5789_3 ( .fault(fault), .net(N5789), .FEN(FEN[2166]), .op(N5789_t3) );
fim FAN_N5789_4 ( .fault(fault), .net(N5789), .FEN(FEN[2167]), .op(N5789_t4) );
fim FAN_N5789_5 ( .fault(fault), .net(N5789), .FEN(FEN[2168]), .op(N5789_t5) );
fim FAN_N5789_6 ( .fault(fault), .net(N5789), .FEN(FEN[2169]), .op(N5789_t6) );
fim FAN_N5789_7 ( .fault(fault), .net(N5789), .FEN(FEN[2170]), .op(N5789_t7) );
fim FAN_N5789_8 ( .fault(fault), .net(N5789), .FEN(FEN[2171]), .op(N5789_t8) );
fim FAN_N5778_0 ( .fault(fault), .net(N5778), .FEN(FEN[2172]), .op(N5778_t0) );
fim FAN_N5778_1 ( .fault(fault), .net(N5778), .FEN(FEN[2173]), .op(N5778_t1) );
fim FAN_N5778_2 ( .fault(fault), .net(N5778), .FEN(FEN[2174]), .op(N5778_t2) );
fim FAN_N5778_3 ( .fault(fault), .net(N5778), .FEN(FEN[2175]), .op(N5778_t3) );
fim FAN_N5778_4 ( .fault(fault), .net(N5778), .FEN(FEN[2176]), .op(N5778_t4) );
fim FAN_N5778_5 ( .fault(fault), .net(N5778), .FEN(FEN[2177]), .op(N5778_t5) );
fim FAN_N5778_6 ( .fault(fault), .net(N5778), .FEN(FEN[2178]), .op(N5778_t6) );
fim FAN_N5778_7 ( .fault(fault), .net(N5778), .FEN(FEN[2179]), .op(N5778_t7) );
fim FAN_N5778_8 ( .fault(fault), .net(N5778), .FEN(FEN[2180]), .op(N5778_t8) );
fim FAN_N5778_9 ( .fault(fault), .net(N5778), .FEN(FEN[2181]), .op(N5778_t9) );
fim FAN_N5771_0 ( .fault(fault), .net(N5771), .FEN(FEN[2182]), .op(N5771_t0) );
fim FAN_N5771_1 ( .fault(fault), .net(N5771), .FEN(FEN[2183]), .op(N5771_t1) );
fim FAN_N5771_2 ( .fault(fault), .net(N5771), .FEN(FEN[2184]), .op(N5771_t2) );
fim FAN_N5771_3 ( .fault(fault), .net(N5771), .FEN(FEN[2185]), .op(N5771_t3) );
fim FAN_N5771_4 ( .fault(fault), .net(N5771), .FEN(FEN[2186]), .op(N5771_t4) );
fim FAN_N5771_5 ( .fault(fault), .net(N5771), .FEN(FEN[2187]), .op(N5771_t5) );
fim FAN_N3169_0 ( .fault(fault), .net(N3169), .FEN(FEN[2188]), .op(N3169_t0) );
fim FAN_N3169_1 ( .fault(fault), .net(N3169), .FEN(FEN[2189]), .op(N3169_t1) );
fim FAN_N3169_2 ( .fault(fault), .net(N3169), .FEN(FEN[2190]), .op(N3169_t2) );
fim FAN_N3173_0 ( .fault(fault), .net(N3173), .FEN(FEN[2191]), .op(N3173_t0) );
fim FAN_N3173_1 ( .fault(fault), .net(N3173), .FEN(FEN[2192]), .op(N3173_t1) );
fim FAN_N3173_2 ( .fault(fault), .net(N3173), .FEN(FEN[2193]), .op(N3173_t2) );
fim FAN_N3173_3 ( .fault(fault), .net(N3173), .FEN(FEN[2194]), .op(N3173_t3) );
fim FAN_N5856_0 ( .fault(fault), .net(N5856), .FEN(FEN[2195]), .op(N5856_t0) );
fim FAN_N5856_1 ( .fault(fault), .net(N5856), .FEN(FEN[2196]), .op(N5856_t1) );
fim FAN_N5856_2 ( .fault(fault), .net(N5856), .FEN(FEN[2197]), .op(N5856_t2) );
fim FAN_N5856_3 ( .fault(fault), .net(N5856), .FEN(FEN[2198]), .op(N5856_t3) );
fim FAN_N5856_4 ( .fault(fault), .net(N5856), .FEN(FEN[2199]), .op(N5856_t4) );
fim FAN_N5856_5 ( .fault(fault), .net(N5856), .FEN(FEN[2200]), .op(N5856_t5) );
fim FAN_N5837_0 ( .fault(fault), .net(N5837), .FEN(FEN[2201]), .op(N5837_t0) );
fim FAN_N5837_1 ( .fault(fault), .net(N5837), .FEN(FEN[2202]), .op(N5837_t1) );
fim FAN_N5837_2 ( .fault(fault), .net(N5837), .FEN(FEN[2203]), .op(N5837_t2) );
fim FAN_N5837_3 ( .fault(fault), .net(N5837), .FEN(FEN[2204]), .op(N5837_t3) );
fim FAN_N5837_4 ( .fault(fault), .net(N5837), .FEN(FEN[2205]), .op(N5837_t4) );
fim FAN_N5837_5 ( .fault(fault), .net(N5837), .FEN(FEN[2206]), .op(N5837_t5) );
fim FAN_N5837_6 ( .fault(fault), .net(N5837), .FEN(FEN[2207]), .op(N5837_t6) );
fim FAN_N5837_7 ( .fault(fault), .net(N5837), .FEN(FEN[2208]), .op(N5837_t7) );
fim FAN_N5837_8 ( .fault(fault), .net(N5837), .FEN(FEN[2209]), .op(N5837_t8) );
fim FAN_N5837_9 ( .fault(fault), .net(N5837), .FEN(FEN[2210]), .op(N5837_t9) );
fim FAN_N5837_10 ( .fault(fault), .net(N5837), .FEN(FEN[2211]), .op(N5837_t10) );
fim FAN_N5837_11 ( .fault(fault), .net(N5837), .FEN(FEN[2212]), .op(N5837_t11) );
fim FAN_N5821_0 ( .fault(fault), .net(N5821), .FEN(FEN[2213]), .op(N5821_t0) );
fim FAN_N5821_1 ( .fault(fault), .net(N5821), .FEN(FEN[2214]), .op(N5821_t1) );
fim FAN_N5821_2 ( .fault(fault), .net(N5821), .FEN(FEN[2215]), .op(N5821_t2) );
fim FAN_N5821_3 ( .fault(fault), .net(N5821), .FEN(FEN[2216]), .op(N5821_t3) );
fim FAN_N5821_4 ( .fault(fault), .net(N5821), .FEN(FEN[2217]), .op(N5821_t4) );
fim FAN_N5821_5 ( .fault(fault), .net(N5821), .FEN(FEN[2218]), .op(N5821_t5) );
fim FAN_N5821_6 ( .fault(fault), .net(N5821), .FEN(FEN[2219]), .op(N5821_t6) );
fim FAN_N5821_7 ( .fault(fault), .net(N5821), .FEN(FEN[2220]), .op(N5821_t7) );
fim FAN_N5821_8 ( .fault(fault), .net(N5821), .FEN(FEN[2221]), .op(N5821_t8) );
fim FAN_N5821_9 ( .fault(fault), .net(N5821), .FEN(FEN[2222]), .op(N5821_t9) );
fim FAN_N5821_10 ( .fault(fault), .net(N5821), .FEN(FEN[2223]), .op(N5821_t10) );
fim FAN_N5821_11 ( .fault(fault), .net(N5821), .FEN(FEN[2224]), .op(N5821_t11) );
fim FAN_N5821_12 ( .fault(fault), .net(N5821), .FEN(FEN[2225]), .op(N5821_t12) );
fim FAN_N5821_13 ( .fault(fault), .net(N5821), .FEN(FEN[2226]), .op(N5821_t13) );
fim FAN_N5821_14 ( .fault(fault), .net(N5821), .FEN(FEN[2227]), .op(N5821_t14) );
fim FAN_N5807_0 ( .fault(fault), .net(N5807), .FEN(FEN[2228]), .op(N5807_t0) );
fim FAN_N5807_1 ( .fault(fault), .net(N5807), .FEN(FEN[2229]), .op(N5807_t1) );
fim FAN_N5807_2 ( .fault(fault), .net(N5807), .FEN(FEN[2230]), .op(N5807_t2) );
fim FAN_N5807_3 ( .fault(fault), .net(N5807), .FEN(FEN[2231]), .op(N5807_t3) );
fim FAN_N5807_4 ( .fault(fault), .net(N5807), .FEN(FEN[2232]), .op(N5807_t4) );
fim FAN_N5807_5 ( .fault(fault), .net(N5807), .FEN(FEN[2233]), .op(N5807_t5) );
fim FAN_N5807_6 ( .fault(fault), .net(N5807), .FEN(FEN[2234]), .op(N5807_t6) );
fim FAN_N5807_7 ( .fault(fault), .net(N5807), .FEN(FEN[2235]), .op(N5807_t7) );
fim FAN_N5807_8 ( .fault(fault), .net(N5807), .FEN(FEN[2236]), .op(N5807_t8) );
fim FAN_N5807_9 ( .fault(fault), .net(N5807), .FEN(FEN[2237]), .op(N5807_t9) );
fim FAN_N5807_10 ( .fault(fault), .net(N5807), .FEN(FEN[2238]), .op(N5807_t10) );
fim FAN_N5807_11 ( .fault(fault), .net(N5807), .FEN(FEN[2239]), .op(N5807_t11) );
fim FAN_N5807_12 ( .fault(fault), .net(N5807), .FEN(FEN[2240]), .op(N5807_t12) );
fim FAN_N5799_0 ( .fault(fault), .net(N5799), .FEN(FEN[2241]), .op(N5799_t0) );
fim FAN_N5799_1 ( .fault(fault), .net(N5799), .FEN(FEN[2242]), .op(N5799_t1) );
fim FAN_N5799_2 ( .fault(fault), .net(N5799), .FEN(FEN[2243]), .op(N5799_t2) );
fim FAN_N5799_3 ( .fault(fault), .net(N5799), .FEN(FEN[2244]), .op(N5799_t3) );
fim FAN_N5799_4 ( .fault(fault), .net(N5799), .FEN(FEN[2245]), .op(N5799_t4) );
fim FAN_N5799_5 ( .fault(fault), .net(N5799), .FEN(FEN[2246]), .op(N5799_t5) );
fim FAN_N5799_6 ( .fault(fault), .net(N5799), .FEN(FEN[2247]), .op(N5799_t6) );
fim FAN_N3185_0 ( .fault(fault), .net(N3185), .FEN(FEN[2248]), .op(N3185_t0) );
fim FAN_N3185_1 ( .fault(fault), .net(N3185), .FEN(FEN[2249]), .op(N3185_t1) );
fim FAN_N3185_2 ( .fault(fault), .net(N3185), .FEN(FEN[2250]), .op(N3185_t2) );
fim FAN_N3189_0 ( .fault(fault), .net(N3189), .FEN(FEN[2251]), .op(N3189_t0) );
fim FAN_N3189_1 ( .fault(fault), .net(N3189), .FEN(FEN[2252]), .op(N3189_t1) );
fim FAN_N3189_2 ( .fault(fault), .net(N3189), .FEN(FEN[2253]), .op(N3189_t2) );
fim FAN_N3189_3 ( .fault(fault), .net(N3189), .FEN(FEN[2254]), .op(N3189_t3) );
fim FAN_N3189_4 ( .fault(fault), .net(N3189), .FEN(FEN[2255]), .op(N3189_t4) );
fim FAN_N3195_0 ( .fault(fault), .net(N3195), .FEN(FEN[2256]), .op(N3195_t0) );
fim FAN_N3195_1 ( .fault(fault), .net(N3195), .FEN(FEN[2257]), .op(N3195_t1) );
fim FAN_N3195_2 ( .fault(fault), .net(N3195), .FEN(FEN[2258]), .op(N3195_t2) );
fim FAN_N3195_3 ( .fault(fault), .net(N3195), .FEN(FEN[2259]), .op(N3195_t3) );
fim FAN_N3195_4 ( .fault(fault), .net(N3195), .FEN(FEN[2260]), .op(N3195_t4) );
fim FAN_N3195_5 ( .fault(fault), .net(N3195), .FEN(FEN[2261]), .op(N3195_t5) );
fim FAN_N5870_0 ( .fault(fault), .net(N5870), .FEN(FEN[2262]), .op(N5870_t0) );
fim FAN_N5870_1 ( .fault(fault), .net(N5870), .FEN(FEN[2263]), .op(N5870_t1) );
fim FAN_N5870_2 ( .fault(fault), .net(N5870), .FEN(FEN[2264]), .op(N5870_t2) );
fim FAN_N5870_3 ( .fault(fault), .net(N5870), .FEN(FEN[2265]), .op(N5870_t3) );
fim FAN_N5870_4 ( .fault(fault), .net(N5870), .FEN(FEN[2266]), .op(N5870_t4) );
fim FAN_N5870_5 ( .fault(fault), .net(N5870), .FEN(FEN[2267]), .op(N5870_t5) );
fim FAN_N5870_6 ( .fault(fault), .net(N5870), .FEN(FEN[2268]), .op(N5870_t6) );
fim FAN_N5870_7 ( .fault(fault), .net(N5870), .FEN(FEN[2269]), .op(N5870_t7) );
fim FAN_N5870_8 ( .fault(fault), .net(N5870), .FEN(FEN[2270]), .op(N5870_t8) );
fim FAN_N5870_9 ( .fault(fault), .net(N5870), .FEN(FEN[2271]), .op(N5870_t9) );
fim FAN_N5881_0 ( .fault(fault), .net(N5881), .FEN(FEN[2272]), .op(N5881_t0) );
fim FAN_N5881_1 ( .fault(fault), .net(N5881), .FEN(FEN[2273]), .op(N5881_t1) );
fim FAN_N5881_2 ( .fault(fault), .net(N5881), .FEN(FEN[2274]), .op(N5881_t2) );
fim FAN_N5881_3 ( .fault(fault), .net(N5881), .FEN(FEN[2275]), .op(N5881_t3) );
fim FAN_N5881_4 ( .fault(fault), .net(N5881), .FEN(FEN[2276]), .op(N5881_t4) );
fim FAN_N5881_5 ( .fault(fault), .net(N5881), .FEN(FEN[2277]), .op(N5881_t5) );
fim FAN_N5881_6 ( .fault(fault), .net(N5881), .FEN(FEN[2278]), .op(N5881_t6) );
fim FAN_N5881_7 ( .fault(fault), .net(N5881), .FEN(FEN[2279]), .op(N5881_t7) );
fim FAN_N5881_8 ( .fault(fault), .net(N5881), .FEN(FEN[2280]), .op(N5881_t8) );
fim FAN_N5881_9 ( .fault(fault), .net(N5881), .FEN(FEN[2281]), .op(N5881_t9) );
fim FAN_N5863_0 ( .fault(fault), .net(N5863), .FEN(FEN[2282]), .op(N5863_t0) );
fim FAN_N5863_1 ( .fault(fault), .net(N5863), .FEN(FEN[2283]), .op(N5863_t1) );
fim FAN_N5863_2 ( .fault(fault), .net(N5863), .FEN(FEN[2284]), .op(N5863_t2) );
fim FAN_N5863_3 ( .fault(fault), .net(N5863), .FEN(FEN[2285]), .op(N5863_t3) );
fim FAN_N5863_4 ( .fault(fault), .net(N5863), .FEN(FEN[2286]), .op(N5863_t4) );
fim FAN_N5863_5 ( .fault(fault), .net(N5863), .FEN(FEN[2287]), .op(N5863_t5) );
fim FAN_N3211_0 ( .fault(fault), .net(N3211), .FEN(FEN[2288]), .op(N3211_t0) );
fim FAN_N3211_1 ( .fault(fault), .net(N3211), .FEN(FEN[2289]), .op(N3211_t1) );
fim FAN_N3211_2 ( .fault(fault), .net(N3211), .FEN(FEN[2290]), .op(N3211_t2) );
fim FAN_N3215_0 ( .fault(fault), .net(N3215), .FEN(FEN[2291]), .op(N3215_t0) );
fim FAN_N3215_1 ( .fault(fault), .net(N3215), .FEN(FEN[2292]), .op(N3215_t1) );
fim FAN_N3215_2 ( .fault(fault), .net(N3215), .FEN(FEN[2293]), .op(N3215_t2) );
fim FAN_N3215_3 ( .fault(fault), .net(N3215), .FEN(FEN[2294]), .op(N3215_t3) );
fim FAN_N3215_4 ( .fault(fault), .net(N3215), .FEN(FEN[2295]), .op(N3215_t4) );
fim FAN_N5905_0 ( .fault(fault), .net(N5905), .FEN(FEN[2296]), .op(N5905_t0) );
fim FAN_N5905_1 ( .fault(fault), .net(N5905), .FEN(FEN[2297]), .op(N5905_t1) );
fim FAN_N5905_2 ( .fault(fault), .net(N5905), .FEN(FEN[2298]), .op(N5905_t2) );
fim FAN_N5905_3 ( .fault(fault), .net(N5905), .FEN(FEN[2299]), .op(N5905_t3) );
fim FAN_N5905_4 ( .fault(fault), .net(N5905), .FEN(FEN[2300]), .op(N5905_t4) );
fim FAN_N5905_5 ( .fault(fault), .net(N5905), .FEN(FEN[2301]), .op(N5905_t5) );
fim FAN_N5905_6 ( .fault(fault), .net(N5905), .FEN(FEN[2302]), .op(N5905_t6) );
fim FAN_N5905_7 ( .fault(fault), .net(N5905), .FEN(FEN[2303]), .op(N5905_t7) );
fim FAN_N5905_8 ( .fault(fault), .net(N5905), .FEN(FEN[2304]), .op(N5905_t8) );
fim FAN_N5936_0 ( .fault(fault), .net(N5936), .FEN(FEN[2305]), .op(N5936_t0) );
fim FAN_N5936_1 ( .fault(fault), .net(N5936), .FEN(FEN[2306]), .op(N5936_t1) );
fim FAN_N5936_2 ( .fault(fault), .net(N5936), .FEN(FEN[2307]), .op(N5936_t2) );
fim FAN_N5936_3 ( .fault(fault), .net(N5936), .FEN(FEN[2308]), .op(N5936_t3) );
fim FAN_N5936_4 ( .fault(fault), .net(N5936), .FEN(FEN[2309]), .op(N5936_t4) );
fim FAN_N5936_5 ( .fault(fault), .net(N5936), .FEN(FEN[2310]), .op(N5936_t5) );
fim FAN_N5915_0 ( .fault(fault), .net(N5915), .FEN(FEN[2311]), .op(N5915_t0) );
fim FAN_N5915_1 ( .fault(fault), .net(N5915), .FEN(FEN[2312]), .op(N5915_t1) );
fim FAN_N5915_2 ( .fault(fault), .net(N5915), .FEN(FEN[2313]), .op(N5915_t2) );
fim FAN_N5915_3 ( .fault(fault), .net(N5915), .FEN(FEN[2314]), .op(N5915_t3) );
fim FAN_N5915_4 ( .fault(fault), .net(N5915), .FEN(FEN[2315]), .op(N5915_t4) );
fim FAN_N5915_5 ( .fault(fault), .net(N5915), .FEN(FEN[2316]), .op(N5915_t5) );
fim FAN_N5915_6 ( .fault(fault), .net(N5915), .FEN(FEN[2317]), .op(N5915_t6) );
fim FAN_N5915_7 ( .fault(fault), .net(N5915), .FEN(FEN[2318]), .op(N5915_t7) );
fim FAN_N5915_8 ( .fault(fault), .net(N5915), .FEN(FEN[2319]), .op(N5915_t8) );
fim FAN_N5915_9 ( .fault(fault), .net(N5915), .FEN(FEN[2320]), .op(N5915_t9) );
fim FAN_N5898_0 ( .fault(fault), .net(N5898), .FEN(FEN[2321]), .op(N5898_t0) );
fim FAN_N5898_1 ( .fault(fault), .net(N5898), .FEN(FEN[2322]), .op(N5898_t1) );
fim FAN_N5898_2 ( .fault(fault), .net(N5898), .FEN(FEN[2323]), .op(N5898_t2) );
fim FAN_N5898_3 ( .fault(fault), .net(N5898), .FEN(FEN[2324]), .op(N5898_t3) );
fim FAN_N5898_4 ( .fault(fault), .net(N5898), .FEN(FEN[2325]), .op(N5898_t4) );
fim FAN_N5898_5 ( .fault(fault), .net(N5898), .FEN(FEN[2326]), .op(N5898_t5) );
fim FAN_N5926_0 ( .fault(fault), .net(N5926), .FEN(FEN[2327]), .op(N5926_t0) );
fim FAN_N5926_1 ( .fault(fault), .net(N5926), .FEN(FEN[2328]), .op(N5926_t1) );
fim FAN_N5926_2 ( .fault(fault), .net(N5926), .FEN(FEN[2329]), .op(N5926_t2) );
fim FAN_N5926_3 ( .fault(fault), .net(N5926), .FEN(FEN[2330]), .op(N5926_t3) );
fim FAN_N5926_4 ( .fault(fault), .net(N5926), .FEN(FEN[2331]), .op(N5926_t4) );
fim FAN_N5926_5 ( .fault(fault), .net(N5926), .FEN(FEN[2332]), .op(N5926_t5) );
fim FAN_N5926_6 ( .fault(fault), .net(N5926), .FEN(FEN[2333]), .op(N5926_t6) );
fim FAN_N5926_7 ( .fault(fault), .net(N5926), .FEN(FEN[2334]), .op(N5926_t7) );
fim FAN_N5926_8 ( .fault(fault), .net(N5926), .FEN(FEN[2335]), .op(N5926_t8) );
fim FAN_N3229_0 ( .fault(fault), .net(N3229), .FEN(FEN[2336]), .op(N3229_t0) );
fim FAN_N3229_1 ( .fault(fault), .net(N3229), .FEN(FEN[2337]), .op(N3229_t1) );
fim FAN_N3232_0 ( .fault(fault), .net(N3232), .FEN(FEN[2338]), .op(N3232_t0) );
fim FAN_N3232_1 ( .fault(fault), .net(N3232), .FEN(FEN[2339]), .op(N3232_t1) );
fim FAN_N3232_2 ( .fault(fault), .net(N3232), .FEN(FEN[2340]), .op(N3232_t2) );
fim FAN_N3236_0 ( .fault(fault), .net(N3236), .FEN(FEN[2341]), .op(N3236_t0) );
fim FAN_N3236_1 ( .fault(fault), .net(N3236), .FEN(FEN[2342]), .op(N3236_t1) );
fim FAN_N3236_2 ( .fault(fault), .net(N3236), .FEN(FEN[2343]), .op(N3236_t2) );
fim FAN_N3236_3 ( .fault(fault), .net(N3236), .FEN(FEN[2344]), .op(N3236_t3) );
fim FAN_N3241_0 ( .fault(fault), .net(N3241), .FEN(FEN[2345]), .op(N3241_t0) );
fim FAN_N3241_1 ( .fault(fault), .net(N3241), .FEN(FEN[2346]), .op(N3241_t1) );
fim FAN_N3241_2 ( .fault(fault), .net(N3241), .FEN(FEN[2347]), .op(N3241_t2) );
fim FAN_N3241_3 ( .fault(fault), .net(N3241), .FEN(FEN[2348]), .op(N3241_t3) );
fim FAN_N3241_4 ( .fault(fault), .net(N3241), .FEN(FEN[2349]), .op(N3241_t4) );
fim FAN_N6204_0 ( .fault(fault), .net(N6204), .FEN(FEN[2350]), .op(N6204_t0) );
fim FAN_N6204_1 ( .fault(fault), .net(N6204), .FEN(FEN[2351]), .op(N6204_t1) );
fim FAN_N6207_0 ( .fault(fault), .net(N6207), .FEN(FEN[2352]), .op(N6207_t0) );
fim FAN_N6207_1 ( .fault(fault), .net(N6207), .FEN(FEN[2353]), .op(N6207_t1) );
fim FAN_N6210_0 ( .fault(fault), .net(N6210), .FEN(FEN[2354]), .op(N6210_t0) );
fim FAN_N6210_1 ( .fault(fault), .net(N6210), .FEN(FEN[2355]), .op(N6210_t1) );
fim FAN_N6000_0 ( .fault(fault), .net(N6000), .FEN(FEN[2356]), .op(N6000_t0) );
fim FAN_N6000_1 ( .fault(fault), .net(N6000), .FEN(FEN[2357]), .op(N6000_t1) );
fim FAN_N5996_0 ( .fault(fault), .net(N5996), .FEN(FEN[2358]), .op(N5996_t0) );
fim FAN_N5996_1 ( .fault(fault), .net(N5996), .FEN(FEN[2359]), .op(N5996_t1) );
fim FAN_N5996_2 ( .fault(fault), .net(N5996), .FEN(FEN[2360]), .op(N5996_t2) );
fim FAN_N5991_0 ( .fault(fault), .net(N5991), .FEN(FEN[2361]), .op(N5991_t0) );
fim FAN_N5991_1 ( .fault(fault), .net(N5991), .FEN(FEN[2362]), .op(N5991_t1) );
fim FAN_N5991_2 ( .fault(fault), .net(N5991), .FEN(FEN[2363]), .op(N5991_t2) );
fim FAN_N5991_3 ( .fault(fault), .net(N5991), .FEN(FEN[2364]), .op(N5991_t3) );
fim FAN_N6018_0 ( .fault(fault), .net(N6018), .FEN(FEN[2365]), .op(N6018_t0) );
fim FAN_N6018_1 ( .fault(fault), .net(N6018), .FEN(FEN[2366]), .op(N6018_t1) );
fim FAN_N6014_0 ( .fault(fault), .net(N6014), .FEN(FEN[2367]), .op(N6014_t0) );
fim FAN_N6014_1 ( .fault(fault), .net(N6014), .FEN(FEN[2368]), .op(N6014_t1) );
fim FAN_N6014_2 ( .fault(fault), .net(N6014), .FEN(FEN[2369]), .op(N6014_t2) );
fim FAN_N6009_0 ( .fault(fault), .net(N6009), .FEN(FEN[2370]), .op(N6009_t0) );
fim FAN_N6009_1 ( .fault(fault), .net(N6009), .FEN(FEN[2371]), .op(N6009_t1) );
fim FAN_N6009_2 ( .fault(fault), .net(N6009), .FEN(FEN[2372]), .op(N6009_t2) );
fim FAN_N6009_3 ( .fault(fault), .net(N6009), .FEN(FEN[2373]), .op(N6009_t3) );
fim FAN_N6003_0 ( .fault(fault), .net(N6003), .FEN(FEN[2374]), .op(N6003_t0) );
fim FAN_N6003_1 ( .fault(fault), .net(N6003), .FEN(FEN[2375]), .op(N6003_t1) );
fim FAN_N6003_2 ( .fault(fault), .net(N6003), .FEN(FEN[2376]), .op(N6003_t2) );
fim FAN_N6003_3 ( .fault(fault), .net(N6003), .FEN(FEN[2377]), .op(N6003_t3) );
fim FAN_N6003_4 ( .fault(fault), .net(N6003), .FEN(FEN[2378]), .op(N6003_t4) );
fim FAN_N6056_0 ( .fault(fault), .net(N6056), .FEN(FEN[2379]), .op(N6056_t0) );
fim FAN_N6056_1 ( .fault(fault), .net(N6056), .FEN(FEN[2380]), .op(N6056_t1) );
fim FAN_N6052_0 ( .fault(fault), .net(N6052), .FEN(FEN[2381]), .op(N6052_t0) );
fim FAN_N6052_1 ( .fault(fault), .net(N6052), .FEN(FEN[2382]), .op(N6052_t1) );
fim FAN_N6052_2 ( .fault(fault), .net(N6052), .FEN(FEN[2383]), .op(N6052_t2) );
fim FAN_N6047_0 ( .fault(fault), .net(N6047), .FEN(FEN[2384]), .op(N6047_t0) );
fim FAN_N6047_1 ( .fault(fault), .net(N6047), .FEN(FEN[2385]), .op(N6047_t1) );
fim FAN_N6047_2 ( .fault(fault), .net(N6047), .FEN(FEN[2386]), .op(N6047_t2) );
fim FAN_N6047_3 ( .fault(fault), .net(N6047), .FEN(FEN[2387]), .op(N6047_t3) );
fim FAN_N6041_0 ( .fault(fault), .net(N6041), .FEN(FEN[2388]), .op(N6041_t0) );
fim FAN_N6041_1 ( .fault(fault), .net(N6041), .FEN(FEN[2389]), .op(N6041_t1) );
fim FAN_N6041_2 ( .fault(fault), .net(N6041), .FEN(FEN[2390]), .op(N6041_t2) );
fim FAN_N6041_3 ( .fault(fault), .net(N6041), .FEN(FEN[2391]), .op(N6041_t3) );
fim FAN_N6041_4 ( .fault(fault), .net(N6041), .FEN(FEN[2392]), .op(N6041_t4) );
fim FAN_N6220_0 ( .fault(fault), .net(N6220), .FEN(FEN[2393]), .op(N6220_t0) );
fim FAN_N6220_1 ( .fault(fault), .net(N6220), .FEN(FEN[2394]), .op(N6220_t1) );
fim FAN_N6079_0 ( .fault(fault), .net(N6079), .FEN(FEN[2395]), .op(N6079_t0) );
fim FAN_N6079_1 ( .fault(fault), .net(N6079), .FEN(FEN[2396]), .op(N6079_t1) );
fim FAN_N6079_2 ( .fault(fault), .net(N6079), .FEN(FEN[2397]), .op(N6079_t2) );
fim FAN_N6083_0 ( .fault(fault), .net(N6083), .FEN(FEN[2398]), .op(N6083_t0) );
fim FAN_N6083_1 ( .fault(fault), .net(N6083), .FEN(FEN[2399]), .op(N6083_t1) );
fim FAN_N6083_2 ( .fault(fault), .net(N6083), .FEN(FEN[2400]), .op(N6083_t2) );
fim FAN_N6087_0 ( .fault(fault), .net(N6087), .FEN(FEN[2401]), .op(N6087_t0) );
fim FAN_N6087_1 ( .fault(fault), .net(N6087), .FEN(FEN[2402]), .op(N6087_t1) );
fim FAN_N6127_0 ( .fault(fault), .net(N6127), .FEN(FEN[2403]), .op(N6127_t0) );
fim FAN_N6127_1 ( .fault(fault), .net(N6127), .FEN(FEN[2404]), .op(N6127_t1) );
fim FAN_N6127_2 ( .fault(fault), .net(N6127), .FEN(FEN[2405]), .op(N6127_t2) );
fim FAN_N6131_0 ( .fault(fault), .net(N6131), .FEN(FEN[2406]), .op(N6131_t0) );
fim FAN_N6131_1 ( .fault(fault), .net(N6131), .FEN(FEN[2407]), .op(N6131_t1) );
fim FAN_N6131_2 ( .fault(fault), .net(N6131), .FEN(FEN[2408]), .op(N6131_t2) );
fim FAN_N6137_0 ( .fault(fault), .net(N6137), .FEN(FEN[2409]), .op(N6137_t0) );
fim FAN_N6137_1 ( .fault(fault), .net(N6137), .FEN(FEN[2410]), .op(N6137_t1) );
fim FAN_N6137_2 ( .fault(fault), .net(N6137), .FEN(FEN[2411]), .op(N6137_t2) );
fim FAN_N6141_0 ( .fault(fault), .net(N6141), .FEN(FEN[2412]), .op(N6141_t0) );
fim FAN_N6141_1 ( .fault(fault), .net(N6141), .FEN(FEN[2413]), .op(N6141_t1) );
fim FAN_N6141_2 ( .fault(fault), .net(N6141), .FEN(FEN[2414]), .op(N6141_t2) );
fim FAN_N6145_0 ( .fault(fault), .net(N6145), .FEN(FEN[2415]), .op(N6145_t0) );
fim FAN_N6145_1 ( .fault(fault), .net(N6145), .FEN(FEN[2416]), .op(N6145_t1) );
fim FAN_N6166_0 ( .fault(fault), .net(N6166), .FEN(FEN[2417]), .op(N6166_t0) );
fim FAN_N6166_1 ( .fault(fault), .net(N6166), .FEN(FEN[2418]), .op(N6166_t1) );
fim FAN_N6166_2 ( .fault(fault), .net(N6166), .FEN(FEN[2419]), .op(N6166_t2) );
fim FAN_N6170_0 ( .fault(fault), .net(N6170), .FEN(FEN[2420]), .op(N6170_t0) );
fim FAN_N6170_1 ( .fault(fault), .net(N6170), .FEN(FEN[2421]), .op(N6170_t1) );
fim FAN_N6170_2 ( .fault(fault), .net(N6170), .FEN(FEN[2422]), .op(N6170_t2) );
fim FAN_N6177_0 ( .fault(fault), .net(N6177), .FEN(FEN[2423]), .op(N6177_t0) );
fim FAN_N6177_1 ( .fault(fault), .net(N6177), .FEN(FEN[2424]), .op(N6177_t1) );
fim FAN_N6177_2 ( .fault(fault), .net(N6177), .FEN(FEN[2425]), .op(N6177_t2) );
fim FAN_N6174_0 ( .fault(fault), .net(N6174), .FEN(FEN[2426]), .op(N6174_t0) );
fim FAN_N6174_1 ( .fault(fault), .net(N6174), .FEN(FEN[2427]), .op(N6174_t1) );
fim FAN_N6196_0 ( .fault(fault), .net(N6196), .FEN(FEN[2428]), .op(N6196_t0) );
fim FAN_N6196_1 ( .fault(fault), .net(N6196), .FEN(FEN[2429]), .op(N6196_t1) );
fim FAN_N6199_0 ( .fault(fault), .net(N6199), .FEN(FEN[2430]), .op(N6199_t0) );
fim FAN_N6199_1 ( .fault(fault), .net(N6199), .FEN(FEN[2431]), .op(N6199_t1) );
fim FAN_N6214_0 ( .fault(fault), .net(N6214), .FEN(FEN[2432]), .op(N6214_t0) );
fim FAN_N6214_1 ( .fault(fault), .net(N6214), .FEN(FEN[2433]), .op(N6214_t1) );
fim FAN_N6217_0 ( .fault(fault), .net(N6217), .FEN(FEN[2434]), .op(N6217_t0) );
fim FAN_N6217_1 ( .fault(fault), .net(N6217), .FEN(FEN[2435]), .op(N6217_t1) );
fim FAN_N5981_0 ( .fault(fault), .net(N5981), .FEN(FEN[2436]), .op(N5981_t0) );
fim FAN_N5981_1 ( .fault(fault), .net(N5981), .FEN(FEN[2437]), .op(N5981_t1) );
fim FAN_N5981_2 ( .fault(fault), .net(N5981), .FEN(FEN[2438]), .op(N5981_t2) );
fim FAN_N5981_3 ( .fault(fault), .net(N5981), .FEN(FEN[2439]), .op(N5981_t3) );
fim FAN_N5981_4 ( .fault(fault), .net(N5981), .FEN(FEN[2440]), .op(N5981_t4) );
fim FAN_N5981_5 ( .fault(fault), .net(N5981), .FEN(FEN[2441]), .op(N5981_t5) );
fim FAN_N5981_6 ( .fault(fault), .net(N5981), .FEN(FEN[2442]), .op(N5981_t6) );
fim FAN_N6249_0 ( .fault(fault), .net(N6249), .FEN(FEN[2443]), .op(N6249_t0) );
fim FAN_N6249_1 ( .fault(fault), .net(N6249), .FEN(FEN[2444]), .op(N6249_t1) );
fim FAN_N6252_0 ( .fault(fault), .net(N6252), .FEN(FEN[2445]), .op(N6252_t0) );
fim FAN_N6252_1 ( .fault(fault), .net(N6252), .FEN(FEN[2446]), .op(N6252_t1) );
fim FAN_N6243_0 ( .fault(fault), .net(N6243), .FEN(FEN[2447]), .op(N6243_t0) );
fim FAN_N6243_1 ( .fault(fault), .net(N6243), .FEN(FEN[2448]), .op(N6243_t1) );
fim FAN_N6246_0 ( .fault(fault), .net(N6246), .FEN(FEN[2449]), .op(N6246_t0) );
fim FAN_N6246_1 ( .fault(fault), .net(N6246), .FEN(FEN[2450]), .op(N6246_t1) );
fim FAN_N6232_0 ( .fault(fault), .net(N6232), .FEN(FEN[2451]), .op(N6232_t0) );
fim FAN_N6232_1 ( .fault(fault), .net(N6232), .FEN(FEN[2452]), .op(N6232_t1) );
fim FAN_N6236_0 ( .fault(fault), .net(N6236), .FEN(FEN[2453]), .op(N6236_t0) );
fim FAN_N6236_1 ( .fault(fault), .net(N6236), .FEN(FEN[2454]), .op(N6236_t1) );
fim FAN_N6263_0 ( .fault(fault), .net(N6263), .FEN(FEN[2455]), .op(N6263_t0) );
fim FAN_N6263_1 ( .fault(fault), .net(N6263), .FEN(FEN[2456]), .op(N6263_t1) );
fim FAN_N6266_0 ( .fault(fault), .net(N6266), .FEN(FEN[2457]), .op(N6266_t0) );
fim FAN_N6266_1 ( .fault(fault), .net(N6266), .FEN(FEN[2458]), .op(N6266_t1) );
fim FAN_N7411_0 ( .fault(fault), .net(N7411), .FEN(FEN[2459]), .op(N7411_t0) );
fim FAN_N7411_1 ( .fault(fault), .net(N7411), .FEN(FEN[2460]), .op(N7411_t1) );
fim FAN_N7414_0 ( .fault(fault), .net(N7414), .FEN(FEN[2461]), .op(N7414_t0) );
fim FAN_N7414_1 ( .fault(fault), .net(N7414), .FEN(FEN[2462]), .op(N7414_t1) );
fim FAN_N7417_0 ( .fault(fault), .net(N7417), .FEN(FEN[2463]), .op(N7417_t0) );
fim FAN_N7417_1 ( .fault(fault), .net(N7417), .FEN(FEN[2464]), .op(N7417_t1) );
fim FAN_N7420_0 ( .fault(fault), .net(N7420), .FEN(FEN[2465]), .op(N7420_t0) );
fim FAN_N7420_1 ( .fault(fault), .net(N7420), .FEN(FEN[2466]), .op(N7420_t1) );
fim FAN_N7423_0 ( .fault(fault), .net(N7423), .FEN(FEN[2467]), .op(N7423_t0) );
fim FAN_N7423_1 ( .fault(fault), .net(N7423), .FEN(FEN[2468]), .op(N7423_t1) );
fim FAN_N7426_0 ( .fault(fault), .net(N7426), .FEN(FEN[2469]), .op(N7426_t0) );
fim FAN_N7426_1 ( .fault(fault), .net(N7426), .FEN(FEN[2470]), .op(N7426_t1) );
fim FAN_N7429_0 ( .fault(fault), .net(N7429), .FEN(FEN[2471]), .op(N7429_t0) );
fim FAN_N7429_1 ( .fault(fault), .net(N7429), .FEN(FEN[2472]), .op(N7429_t1) );
fim FAN_N7432_0 ( .fault(fault), .net(N7432), .FEN(FEN[2473]), .op(N7432_t0) );
fim FAN_N7432_1 ( .fault(fault), .net(N7432), .FEN(FEN[2474]), .op(N7432_t1) );
fim FAN_N7435_0 ( .fault(fault), .net(N7435), .FEN(FEN[2475]), .op(N7435_t0) );
fim FAN_N7435_1 ( .fault(fault), .net(N7435), .FEN(FEN[2476]), .op(N7435_t1) );
fim FAN_N7438_0 ( .fault(fault), .net(N7438), .FEN(FEN[2477]), .op(N7438_t0) );
fim FAN_N7438_1 ( .fault(fault), .net(N7438), .FEN(FEN[2478]), .op(N7438_t1) );
fim FAN_N7136_0 ( .fault(fault), .net(N7136), .FEN(FEN[2479]), .op(N7136_t0) );
fim FAN_N7136_1 ( .fault(fault), .net(N7136), .FEN(FEN[2480]), .op(N7136_t1) );
fim FAN_N7136_2 ( .fault(fault), .net(N7136), .FEN(FEN[2481]), .op(N7136_t2) );
fim FAN_N7136_3 ( .fault(fault), .net(N7136), .FEN(FEN[2482]), .op(N7136_t3) );
fim FAN_N7136_4 ( .fault(fault), .net(N7136), .FEN(FEN[2483]), .op(N7136_t4) );
fim FAN_N6923_0 ( .fault(fault), .net(N6923), .FEN(FEN[2484]), .op(N6923_t0) );
fim FAN_N6923_1 ( .fault(fault), .net(N6923), .FEN(FEN[2485]), .op(N6923_t1) );
fim FAN_N6923_2 ( .fault(fault), .net(N6923), .FEN(FEN[2486]), .op(N6923_t2) );
fim FAN_N6923_3 ( .fault(fault), .net(N6923), .FEN(FEN[2487]), .op(N6923_t3) );
fim FAN_N6923_4 ( .fault(fault), .net(N6923), .FEN(FEN[2488]), .op(N6923_t4) );
fim FAN_N6762_0 ( .fault(fault), .net(N6762), .FEN(FEN[2489]), .op(N6762_t0) );
fim FAN_N6762_1 ( .fault(fault), .net(N6762), .FEN(FEN[2490]), .op(N6762_t1) );
fim FAN_N6762_2 ( .fault(fault), .net(N6762), .FEN(FEN[2491]), .op(N6762_t2) );
fim FAN_N7459_0 ( .fault(fault), .net(N7459), .FEN(FEN[2492]), .op(N7459_t0) );
fim FAN_N7459_1 ( .fault(fault), .net(N7459), .FEN(FEN[2493]), .op(N7459_t1) );
fim FAN_N7462_0 ( .fault(fault), .net(N7462), .FEN(FEN[2494]), .op(N7462_t0) );
fim FAN_N7462_1 ( .fault(fault), .net(N7462), .FEN(FEN[2495]), .op(N7462_t1) );
fim FAN_N6784_0 ( .fault(fault), .net(N6784), .FEN(FEN[2496]), .op(N6784_t0) );
fim FAN_N6784_1 ( .fault(fault), .net(N6784), .FEN(FEN[2497]), .op(N6784_t1) );
fim FAN_N6815_0 ( .fault(fault), .net(N6815), .FEN(FEN[2498]), .op(N6815_t0) );
fim FAN_N6815_1 ( .fault(fault), .net(N6815), .FEN(FEN[2499]), .op(N6815_t1) );
fim FAN_N6818_0 ( .fault(fault), .net(N6818), .FEN(FEN[2500]), .op(N6818_t0) );
fim FAN_N6818_1 ( .fault(fault), .net(N6818), .FEN(FEN[2501]), .op(N6818_t1) );
fim FAN_N6821_0 ( .fault(fault), .net(N6821), .FEN(FEN[2502]), .op(N6821_t0) );
fim FAN_N6821_1 ( .fault(fault), .net(N6821), .FEN(FEN[2503]), .op(N6821_t1) );
fim FAN_N6824_0 ( .fault(fault), .net(N6824), .FEN(FEN[2504]), .op(N6824_t0) );
fim FAN_N6824_1 ( .fault(fault), .net(N6824), .FEN(FEN[2505]), .op(N6824_t1) );
fim FAN_N6827_0 ( .fault(fault), .net(N6827), .FEN(FEN[2506]), .op(N6827_t0) );
fim FAN_N6827_1 ( .fault(fault), .net(N6827), .FEN(FEN[2507]), .op(N6827_t1) );
fim FAN_N6830_0 ( .fault(fault), .net(N6830), .FEN(FEN[2508]), .op(N6830_t0) );
fim FAN_N6830_1 ( .fault(fault), .net(N6830), .FEN(FEN[2509]), .op(N6830_t1) );
fim FAN_N6800_0 ( .fault(fault), .net(N6800), .FEN(FEN[2510]), .op(N6800_t0) );
fim FAN_N6800_1 ( .fault(fault), .net(N6800), .FEN(FEN[2511]), .op(N6800_t1) );
fim FAN_N6797_0 ( .fault(fault), .net(N6797), .FEN(FEN[2512]), .op(N6797_t0) );
fim FAN_N6797_1 ( .fault(fault), .net(N6797), .FEN(FEN[2513]), .op(N6797_t1) );
fim FAN_N6806_0 ( .fault(fault), .net(N6806), .FEN(FEN[2514]), .op(N6806_t0) );
fim FAN_N6806_1 ( .fault(fault), .net(N6806), .FEN(FEN[2515]), .op(N6806_t1) );
fim FAN_N6803_0 ( .fault(fault), .net(N6803), .FEN(FEN[2516]), .op(N6803_t0) );
fim FAN_N6803_1 ( .fault(fault), .net(N6803), .FEN(FEN[2517]), .op(N6803_t1) );
fim FAN_N6812_0 ( .fault(fault), .net(N6812), .FEN(FEN[2518]), .op(N6812_t0) );
fim FAN_N6812_1 ( .fault(fault), .net(N6812), .FEN(FEN[2519]), .op(N6812_t1) );
fim FAN_N6809_0 ( .fault(fault), .net(N6809), .FEN(FEN[2520]), .op(N6809_t0) );
fim FAN_N6809_1 ( .fault(fault), .net(N6809), .FEN(FEN[2521]), .op(N6809_t1) );
fim FAN_N6845_0 ( .fault(fault), .net(N6845), .FEN(FEN[2522]), .op(N6845_t0) );
fim FAN_N6845_1 ( .fault(fault), .net(N6845), .FEN(FEN[2523]), .op(N6845_t1) );
fim FAN_N7488_0 ( .fault(fault), .net(N7488), .FEN(FEN[2524]), .op(N7488_t0) );
fim FAN_N7488_1 ( .fault(fault), .net(N7488), .FEN(FEN[2525]), .op(N7488_t1) );
fim FAN_N7500_0 ( .fault(fault), .net(N7500), .FEN(FEN[2526]), .op(N7500_t0) );
fim FAN_N7500_1 ( .fault(fault), .net(N7500), .FEN(FEN[2527]), .op(N7500_t1) );
fim FAN_N7515_0 ( .fault(fault), .net(N7515), .FEN(FEN[2528]), .op(N7515_t0) );
fim FAN_N7515_1 ( .fault(fault), .net(N7515), .FEN(FEN[2529]), .op(N7515_t1) );
fim FAN_N7518_0 ( .fault(fault), .net(N7518), .FEN(FEN[2530]), .op(N7518_t0) );
fim FAN_N7518_1 ( .fault(fault), .net(N7518), .FEN(FEN[2531]), .op(N7518_t1) );
fim FAN_N6833_0 ( .fault(fault), .net(N6833), .FEN(FEN[2532]), .op(N6833_t0) );
fim FAN_N6833_1 ( .fault(fault), .net(N6833), .FEN(FEN[2533]), .op(N6833_t1) );
fim FAN_N6867_0 ( .fault(fault), .net(N6867), .FEN(FEN[2534]), .op(N6867_t0) );
fim FAN_N6867_1 ( .fault(fault), .net(N6867), .FEN(FEN[2535]), .op(N6867_t1) );
fim FAN_N6881_0 ( .fault(fault), .net(N6881), .FEN(FEN[2536]), .op(N6881_t0) );
fim FAN_N6881_1 ( .fault(fault), .net(N6881), .FEN(FEN[2537]), .op(N6881_t1) );
fim FAN_N7533_0 ( .fault(fault), .net(N7533), .FEN(FEN[2538]), .op(N7533_t0) );
fim FAN_N7533_1 ( .fault(fault), .net(N7533), .FEN(FEN[2539]), .op(N7533_t1) );
fim FAN_N7536_0 ( .fault(fault), .net(N7536), .FEN(FEN[2540]), .op(N7536_t0) );
fim FAN_N7536_1 ( .fault(fault), .net(N7536), .FEN(FEN[2541]), .op(N7536_t1) );
fim FAN_N7539_0 ( .fault(fault), .net(N7539), .FEN(FEN[2542]), .op(N7539_t0) );
fim FAN_N7539_1 ( .fault(fault), .net(N7539), .FEN(FEN[2543]), .op(N7539_t1) );
fim FAN_N7542_0 ( .fault(fault), .net(N7542), .FEN(FEN[2544]), .op(N7542_t0) );
fim FAN_N7542_1 ( .fault(fault), .net(N7542), .FEN(FEN[2545]), .op(N7542_t1) );
fim FAN_N7545_0 ( .fault(fault), .net(N7545), .FEN(FEN[2546]), .op(N7545_t0) );
fim FAN_N7545_1 ( .fault(fault), .net(N7545), .FEN(FEN[2547]), .op(N7545_t1) );
fim FAN_N7548_0 ( .fault(fault), .net(N7548), .FEN(FEN[2548]), .op(N7548_t0) );
fim FAN_N7548_1 ( .fault(fault), .net(N7548), .FEN(FEN[2549]), .op(N7548_t1) );
fim FAN_N6901_0 ( .fault(fault), .net(N6901), .FEN(FEN[2550]), .op(N6901_t0) );
fim FAN_N6901_1 ( .fault(fault), .net(N6901), .FEN(FEN[2551]), .op(N6901_t1) );
fim FAN_N6901_2 ( .fault(fault), .net(N6901), .FEN(FEN[2552]), .op(N6901_t2) );
fim FAN_N6901_3 ( .fault(fault), .net(N6901), .FEN(FEN[2553]), .op(N6901_t3) );
fim FAN_N6901_4 ( .fault(fault), .net(N6901), .FEN(FEN[2554]), .op(N6901_t4) );
fim FAN_N6901_5 ( .fault(fault), .net(N6901), .FEN(FEN[2555]), .op(N6901_t5) );
fim FAN_N6901_6 ( .fault(fault), .net(N6901), .FEN(FEN[2556]), .op(N6901_t6) );
fim FAN_N6901_7 ( .fault(fault), .net(N6901), .FEN(FEN[2557]), .op(N6901_t7) );
fim FAN_N6901_8 ( .fault(fault), .net(N6901), .FEN(FEN[2558]), .op(N6901_t8) );
fim FAN_N6901_9 ( .fault(fault), .net(N6901), .FEN(FEN[2559]), .op(N6901_t9) );
fim FAN_N6912_0 ( .fault(fault), .net(N6912), .FEN(FEN[2560]), .op(N6912_t0) );
fim FAN_N6912_1 ( .fault(fault), .net(N6912), .FEN(FEN[2561]), .op(N6912_t1) );
fim FAN_N6912_2 ( .fault(fault), .net(N6912), .FEN(FEN[2562]), .op(N6912_t2) );
fim FAN_N6912_3 ( .fault(fault), .net(N6912), .FEN(FEN[2563]), .op(N6912_t3) );
fim FAN_N6912_4 ( .fault(fault), .net(N6912), .FEN(FEN[2564]), .op(N6912_t4) );
fim FAN_N6912_5 ( .fault(fault), .net(N6912), .FEN(FEN[2565]), .op(N6912_t5) );
fim FAN_N6912_6 ( .fault(fault), .net(N6912), .FEN(FEN[2566]), .op(N6912_t6) );
fim FAN_N6912_7 ( .fault(fault), .net(N6912), .FEN(FEN[2567]), .op(N6912_t7) );
fim FAN_N6912_8 ( .fault(fault), .net(N6912), .FEN(FEN[2568]), .op(N6912_t8) );
fim FAN_N6912_9 ( .fault(fault), .net(N6912), .FEN(FEN[2569]), .op(N6912_t9) );
fim FAN_N6894_0 ( .fault(fault), .net(N6894), .FEN(FEN[2570]), .op(N6894_t0) );
fim FAN_N6894_1 ( .fault(fault), .net(N6894), .FEN(FEN[2571]), .op(N6894_t1) );
fim FAN_N6894_2 ( .fault(fault), .net(N6894), .FEN(FEN[2572]), .op(N6894_t2) );
fim FAN_N6894_3 ( .fault(fault), .net(N6894), .FEN(FEN[2573]), .op(N6894_t3) );
fim FAN_N6894_4 ( .fault(fault), .net(N6894), .FEN(FEN[2574]), .op(N6894_t4) );
fim FAN_N6894_5 ( .fault(fault), .net(N6894), .FEN(FEN[2575]), .op(N6894_t5) );
fim FAN_N4545_0 ( .fault(fault), .net(N4545), .FEN(FEN[2576]), .op(N4545_t0) );
fim FAN_N4545_1 ( .fault(fault), .net(N4545), .FEN(FEN[2577]), .op(N4545_t1) );
fim FAN_N4545_2 ( .fault(fault), .net(N4545), .FEN(FEN[2578]), .op(N4545_t2) );
fim FAN_N4549_0 ( .fault(fault), .net(N4549), .FEN(FEN[2579]), .op(N4549_t0) );
fim FAN_N4549_1 ( .fault(fault), .net(N4549), .FEN(FEN[2580]), .op(N4549_t1) );
fim FAN_N4549_2 ( .fault(fault), .net(N4549), .FEN(FEN[2581]), .op(N4549_t2) );
fim FAN_N4549_3 ( .fault(fault), .net(N4549), .FEN(FEN[2582]), .op(N4549_t3) );
fim FAN_N4549_4 ( .fault(fault), .net(N4549), .FEN(FEN[2583]), .op(N4549_t4) );
fim FAN_N6929_0 ( .fault(fault), .net(N6929), .FEN(FEN[2584]), .op(N6929_t0) );
fim FAN_N6929_1 ( .fault(fault), .net(N6929), .FEN(FEN[2585]), .op(N6929_t1) );
fim FAN_N6929_2 ( .fault(fault), .net(N6929), .FEN(FEN[2586]), .op(N6929_t2) );
fim FAN_N6929_3 ( .fault(fault), .net(N6929), .FEN(FEN[2587]), .op(N6929_t3) );
fim FAN_N6929_4 ( .fault(fault), .net(N6929), .FEN(FEN[2588]), .op(N6929_t4) );
fim FAN_N6929_5 ( .fault(fault), .net(N6929), .FEN(FEN[2589]), .op(N6929_t5) );
fim FAN_N4563_0 ( .fault(fault), .net(N4563), .FEN(FEN[2590]), .op(N4563_t0) );
fim FAN_N4563_1 ( .fault(fault), .net(N4563), .FEN(FEN[2591]), .op(N4563_t1) );
fim FAN_N6936_0 ( .fault(fault), .net(N6936), .FEN(FEN[2592]), .op(N6936_t0) );
fim FAN_N6936_1 ( .fault(fault), .net(N6936), .FEN(FEN[2593]), .op(N6936_t1) );
fim FAN_N6936_2 ( .fault(fault), .net(N6936), .FEN(FEN[2594]), .op(N6936_t2) );
fim FAN_N6936_3 ( .fault(fault), .net(N6936), .FEN(FEN[2595]), .op(N6936_t3) );
fim FAN_N6936_4 ( .fault(fault), .net(N6936), .FEN(FEN[2596]), .op(N6936_t4) );
fim FAN_N6936_5 ( .fault(fault), .net(N6936), .FEN(FEN[2597]), .op(N6936_t5) );
fim FAN_N6936_6 ( .fault(fault), .net(N6936), .FEN(FEN[2598]), .op(N6936_t6) );
fim FAN_N6936_7 ( .fault(fault), .net(N6936), .FEN(FEN[2599]), .op(N6936_t7) );
fim FAN_N6936_8 ( .fault(fault), .net(N6936), .FEN(FEN[2600]), .op(N6936_t8) );
fim FAN_N4566_0 ( .fault(fault), .net(N4566), .FEN(FEN[2601]), .op(N4566_t0) );
fim FAN_N4566_1 ( .fault(fault), .net(N4566), .FEN(FEN[2602]), .op(N4566_t1) );
fim FAN_N4566_2 ( .fault(fault), .net(N4566), .FEN(FEN[2603]), .op(N4566_t2) );
fim FAN_N6946_0 ( .fault(fault), .net(N6946), .FEN(FEN[2604]), .op(N6946_t0) );
fim FAN_N6946_1 ( .fault(fault), .net(N6946), .FEN(FEN[2605]), .op(N6946_t1) );
fim FAN_N6946_2 ( .fault(fault), .net(N6946), .FEN(FEN[2606]), .op(N6946_t2) );
fim FAN_N6946_3 ( .fault(fault), .net(N6946), .FEN(FEN[2607]), .op(N6946_t3) );
fim FAN_N6946_4 ( .fault(fault), .net(N6946), .FEN(FEN[2608]), .op(N6946_t4) );
fim FAN_N6946_5 ( .fault(fault), .net(N6946), .FEN(FEN[2609]), .op(N6946_t5) );
fim FAN_N6946_6 ( .fault(fault), .net(N6946), .FEN(FEN[2610]), .op(N6946_t6) );
fim FAN_N6946_7 ( .fault(fault), .net(N6946), .FEN(FEN[2611]), .op(N6946_t7) );
fim FAN_N6946_8 ( .fault(fault), .net(N6946), .FEN(FEN[2612]), .op(N6946_t8) );
fim FAN_N6946_9 ( .fault(fault), .net(N6946), .FEN(FEN[2613]), .op(N6946_t9) );
fim FAN_N4570_0 ( .fault(fault), .net(N4570), .FEN(FEN[2614]), .op(N4570_t0) );
fim FAN_N4570_1 ( .fault(fault), .net(N4570), .FEN(FEN[2615]), .op(N4570_t1) );
fim FAN_N4570_2 ( .fault(fault), .net(N4570), .FEN(FEN[2616]), .op(N4570_t2) );
fim FAN_N4570_3 ( .fault(fault), .net(N4570), .FEN(FEN[2617]), .op(N4570_t3) );
fim FAN_N6957_0 ( .fault(fault), .net(N6957), .FEN(FEN[2618]), .op(N6957_t0) );
fim FAN_N6957_1 ( .fault(fault), .net(N6957), .FEN(FEN[2619]), .op(N6957_t1) );
fim FAN_N6957_2 ( .fault(fault), .net(N6957), .FEN(FEN[2620]), .op(N6957_t2) );
fim FAN_N6957_3 ( .fault(fault), .net(N6957), .FEN(FEN[2621]), .op(N6957_t3) );
fim FAN_N6957_4 ( .fault(fault), .net(N6957), .FEN(FEN[2622]), .op(N6957_t4) );
fim FAN_N6957_5 ( .fault(fault), .net(N6957), .FEN(FEN[2623]), .op(N6957_t5) );
fim FAN_N6957_6 ( .fault(fault), .net(N6957), .FEN(FEN[2624]), .op(N6957_t6) );
fim FAN_N6957_7 ( .fault(fault), .net(N6957), .FEN(FEN[2625]), .op(N6957_t7) );
fim FAN_N6957_8 ( .fault(fault), .net(N6957), .FEN(FEN[2626]), .op(N6957_t8) );
fim FAN_N5960_0 ( .fault(fault), .net(N5960), .FEN(FEN[2627]), .op(N5960_t0) );
fim FAN_N5960_1 ( .fault(fault), .net(N5960), .FEN(FEN[2628]), .op(N5960_t1) );
fim FAN_N5960_2 ( .fault(fault), .net(N5960), .FEN(FEN[2629]), .op(N5960_t2) );
fim FAN_N5960_3 ( .fault(fault), .net(N5960), .FEN(FEN[2630]), .op(N5960_t3) );
fim FAN_N5960_4 ( .fault(fault), .net(N5960), .FEN(FEN[2631]), .op(N5960_t4) );
fim FAN_N7049_0 ( .fault(fault), .net(N7049), .FEN(FEN[2632]), .op(N7049_t0) );
fim FAN_N7049_1 ( .fault(fault), .net(N7049), .FEN(FEN[2633]), .op(N7049_t1) );
fim FAN_N7049_2 ( .fault(fault), .net(N7049), .FEN(FEN[2634]), .op(N7049_t2) );
fim FAN_N7049_3 ( .fault(fault), .net(N7049), .FEN(FEN[2635]), .op(N7049_t3) );
fim FAN_N7049_4 ( .fault(fault), .net(N7049), .FEN(FEN[2636]), .op(N7049_t4) );
fim FAN_N6988_0 ( .fault(fault), .net(N6988), .FEN(FEN[2637]), .op(N6988_t0) );
fim FAN_N6988_1 ( .fault(fault), .net(N6988), .FEN(FEN[2638]), .op(N6988_t1) );
fim FAN_N6988_2 ( .fault(fault), .net(N6988), .FEN(FEN[2639]), .op(N6988_t2) );
fim FAN_N6988_3 ( .fault(fault), .net(N6988), .FEN(FEN[2640]), .op(N6988_t3) );
fim FAN_N6988_4 ( .fault(fault), .net(N6988), .FEN(FEN[2641]), .op(N6988_t4) );
fim FAN_N6988_5 ( .fault(fault), .net(N6988), .FEN(FEN[2642]), .op(N6988_t5) );
fim FAN_N6988_6 ( .fault(fault), .net(N6988), .FEN(FEN[2643]), .op(N6988_t6) );
fim FAN_N6988_7 ( .fault(fault), .net(N6988), .FEN(FEN[2644]), .op(N6988_t7) );
fim FAN_N6988_8 ( .fault(fault), .net(N6988), .FEN(FEN[2645]), .op(N6988_t8) );
fim FAN_N6977_0 ( .fault(fault), .net(N6977), .FEN(FEN[2646]), .op(N6977_t0) );
fim FAN_N6977_1 ( .fault(fault), .net(N6977), .FEN(FEN[2647]), .op(N6977_t1) );
fim FAN_N6977_2 ( .fault(fault), .net(N6977), .FEN(FEN[2648]), .op(N6977_t2) );
fim FAN_N6977_3 ( .fault(fault), .net(N6977), .FEN(FEN[2649]), .op(N6977_t3) );
fim FAN_N6977_4 ( .fault(fault), .net(N6977), .FEN(FEN[2650]), .op(N6977_t4) );
fim FAN_N6977_5 ( .fault(fault), .net(N6977), .FEN(FEN[2651]), .op(N6977_t5) );
fim FAN_N6977_6 ( .fault(fault), .net(N6977), .FEN(FEN[2652]), .op(N6977_t6) );
fim FAN_N6977_7 ( .fault(fault), .net(N6977), .FEN(FEN[2653]), .op(N6977_t7) );
fim FAN_N6977_8 ( .fault(fault), .net(N6977), .FEN(FEN[2654]), .op(N6977_t8) );
fim FAN_N6977_9 ( .fault(fault), .net(N6977), .FEN(FEN[2655]), .op(N6977_t9) );
fim FAN_N6970_0 ( .fault(fault), .net(N6970), .FEN(FEN[2656]), .op(N6970_t0) );
fim FAN_N6970_1 ( .fault(fault), .net(N6970), .FEN(FEN[2657]), .op(N6970_t1) );
fim FAN_N6970_2 ( .fault(fault), .net(N6970), .FEN(FEN[2658]), .op(N6970_t2) );
fim FAN_N6970_3 ( .fault(fault), .net(N6970), .FEN(FEN[2659]), .op(N6970_t3) );
fim FAN_N6970_4 ( .fault(fault), .net(N6970), .FEN(FEN[2660]), .op(N6970_t4) );
fim FAN_N6970_5 ( .fault(fault), .net(N6970), .FEN(FEN[2661]), .op(N6970_t5) );
fim FAN_N4577_0 ( .fault(fault), .net(N4577), .FEN(FEN[2662]), .op(N4577_t0) );
fim FAN_N4577_1 ( .fault(fault), .net(N4577), .FEN(FEN[2663]), .op(N4577_t1) );
fim FAN_N4577_2 ( .fault(fault), .net(N4577), .FEN(FEN[2664]), .op(N4577_t2) );
fim FAN_N4581_0 ( .fault(fault), .net(N4581), .FEN(FEN[2665]), .op(N4581_t0) );
fim FAN_N4581_1 ( .fault(fault), .net(N4581), .FEN(FEN[2666]), .op(N4581_t1) );
fim FAN_N4581_2 ( .fault(fault), .net(N4581), .FEN(FEN[2667]), .op(N4581_t2) );
fim FAN_N4581_3 ( .fault(fault), .net(N4581), .FEN(FEN[2668]), .op(N4581_t3) );
fim FAN_N6998_0 ( .fault(fault), .net(N6998), .FEN(FEN[2669]), .op(N6998_t0) );
fim FAN_N6998_1 ( .fault(fault), .net(N6998), .FEN(FEN[2670]), .op(N6998_t1) );
fim FAN_N6998_2 ( .fault(fault), .net(N6998), .FEN(FEN[2671]), .op(N6998_t2) );
fim FAN_N6998_3 ( .fault(fault), .net(N6998), .FEN(FEN[2672]), .op(N6998_t3) );
fim FAN_N6998_4 ( .fault(fault), .net(N6998), .FEN(FEN[2673]), .op(N6998_t4) );
fim FAN_N6998_5 ( .fault(fault), .net(N6998), .FEN(FEN[2674]), .op(N6998_t5) );
fim FAN_N6998_6 ( .fault(fault), .net(N6998), .FEN(FEN[2675]), .op(N6998_t6) );
fim FAN_N4593_0 ( .fault(fault), .net(N4593), .FEN(FEN[2676]), .op(N4593_t0) );
fim FAN_N4593_1 ( .fault(fault), .net(N4593), .FEN(FEN[2677]), .op(N4593_t1) );
fim FAN_N4593_2 ( .fault(fault), .net(N4593), .FEN(FEN[2678]), .op(N4593_t2) );
fim FAN_N7006_0 ( .fault(fault), .net(N7006), .FEN(FEN[2679]), .op(N7006_t0) );
fim FAN_N7006_1 ( .fault(fault), .net(N7006), .FEN(FEN[2680]), .op(N7006_t1) );
fim FAN_N7006_2 ( .fault(fault), .net(N7006), .FEN(FEN[2681]), .op(N7006_t2) );
fim FAN_N7006_3 ( .fault(fault), .net(N7006), .FEN(FEN[2682]), .op(N7006_t3) );
fim FAN_N7006_4 ( .fault(fault), .net(N7006), .FEN(FEN[2683]), .op(N7006_t4) );
fim FAN_N7006_5 ( .fault(fault), .net(N7006), .FEN(FEN[2684]), .op(N7006_t5) );
fim FAN_N7006_6 ( .fault(fault), .net(N7006), .FEN(FEN[2685]), .op(N7006_t6) );
fim FAN_N7006_7 ( .fault(fault), .net(N7006), .FEN(FEN[2686]), .op(N7006_t7) );
fim FAN_N7006_8 ( .fault(fault), .net(N7006), .FEN(FEN[2687]), .op(N7006_t8) );
fim FAN_N7006_9 ( .fault(fault), .net(N7006), .FEN(FEN[2688]), .op(N7006_t9) );
fim FAN_N7006_10 ( .fault(fault), .net(N7006), .FEN(FEN[2689]), .op(N7006_t10) );
fim FAN_N7006_11 ( .fault(fault), .net(N7006), .FEN(FEN[2690]), .op(N7006_t11) );
fim FAN_N7006_12 ( .fault(fault), .net(N7006), .FEN(FEN[2691]), .op(N7006_t12) );
fim FAN_N4597_0 ( .fault(fault), .net(N4597), .FEN(FEN[2692]), .op(N4597_t0) );
fim FAN_N4597_1 ( .fault(fault), .net(N4597), .FEN(FEN[2693]), .op(N4597_t1) );
fim FAN_N4597_2 ( .fault(fault), .net(N4597), .FEN(FEN[2694]), .op(N4597_t2) );
fim FAN_N4597_3 ( .fault(fault), .net(N4597), .FEN(FEN[2695]), .op(N4597_t3) );
fim FAN_N4597_4 ( .fault(fault), .net(N4597), .FEN(FEN[2696]), .op(N4597_t4) );
fim FAN_N7020_0 ( .fault(fault), .net(N7020), .FEN(FEN[2697]), .op(N7020_t0) );
fim FAN_N7020_1 ( .fault(fault), .net(N7020), .FEN(FEN[2698]), .op(N7020_t1) );
fim FAN_N7020_2 ( .fault(fault), .net(N7020), .FEN(FEN[2699]), .op(N7020_t2) );
fim FAN_N7020_3 ( .fault(fault), .net(N7020), .FEN(FEN[2700]), .op(N7020_t3) );
fim FAN_N7020_4 ( .fault(fault), .net(N7020), .FEN(FEN[2701]), .op(N7020_t4) );
fim FAN_N7020_5 ( .fault(fault), .net(N7020), .FEN(FEN[2702]), .op(N7020_t5) );
fim FAN_N7020_6 ( .fault(fault), .net(N7020), .FEN(FEN[2703]), .op(N7020_t6) );
fim FAN_N7020_7 ( .fault(fault), .net(N7020), .FEN(FEN[2704]), .op(N7020_t7) );
fim FAN_N7020_8 ( .fault(fault), .net(N7020), .FEN(FEN[2705]), .op(N7020_t8) );
fim FAN_N7020_9 ( .fault(fault), .net(N7020), .FEN(FEN[2706]), .op(N7020_t9) );
fim FAN_N7020_10 ( .fault(fault), .net(N7020), .FEN(FEN[2707]), .op(N7020_t10) );
fim FAN_N7020_11 ( .fault(fault), .net(N7020), .FEN(FEN[2708]), .op(N7020_t11) );
fim FAN_N7020_12 ( .fault(fault), .net(N7020), .FEN(FEN[2709]), .op(N7020_t12) );
fim FAN_N7020_13 ( .fault(fault), .net(N7020), .FEN(FEN[2710]), .op(N7020_t13) );
fim FAN_N7020_14 ( .fault(fault), .net(N7020), .FEN(FEN[2711]), .op(N7020_t14) );
fim FAN_N4603_0 ( .fault(fault), .net(N4603), .FEN(FEN[2712]), .op(N4603_t0) );
fim FAN_N4603_1 ( .fault(fault), .net(N4603), .FEN(FEN[2713]), .op(N4603_t1) );
fim FAN_N4603_2 ( .fault(fault), .net(N4603), .FEN(FEN[2714]), .op(N4603_t2) );
fim FAN_N4603_3 ( .fault(fault), .net(N4603), .FEN(FEN[2715]), .op(N4603_t3) );
fim FAN_N4603_4 ( .fault(fault), .net(N4603), .FEN(FEN[2716]), .op(N4603_t4) );
fim FAN_N4603_5 ( .fault(fault), .net(N4603), .FEN(FEN[2717]), .op(N4603_t5) );
fim FAN_N7036_0 ( .fault(fault), .net(N7036), .FEN(FEN[2718]), .op(N7036_t0) );
fim FAN_N7036_1 ( .fault(fault), .net(N7036), .FEN(FEN[2719]), .op(N7036_t1) );
fim FAN_N7036_2 ( .fault(fault), .net(N7036), .FEN(FEN[2720]), .op(N7036_t2) );
fim FAN_N7036_3 ( .fault(fault), .net(N7036), .FEN(FEN[2721]), .op(N7036_t3) );
fim FAN_N7036_4 ( .fault(fault), .net(N7036), .FEN(FEN[2722]), .op(N7036_t4) );
fim FAN_N7036_5 ( .fault(fault), .net(N7036), .FEN(FEN[2723]), .op(N7036_t5) );
fim FAN_N7036_6 ( .fault(fault), .net(N7036), .FEN(FEN[2724]), .op(N7036_t6) );
fim FAN_N7036_7 ( .fault(fault), .net(N7036), .FEN(FEN[2725]), .op(N7036_t7) );
fim FAN_N7036_8 ( .fault(fault), .net(N7036), .FEN(FEN[2726]), .op(N7036_t8) );
fim FAN_N7036_9 ( .fault(fault), .net(N7036), .FEN(FEN[2727]), .op(N7036_t9) );
fim FAN_N7036_10 ( .fault(fault), .net(N7036), .FEN(FEN[2728]), .op(N7036_t10) );
fim FAN_N7036_11 ( .fault(fault), .net(N7036), .FEN(FEN[2729]), .op(N7036_t11) );
fim FAN_N7057_0 ( .fault(fault), .net(N7057), .FEN(FEN[2730]), .op(N7057_t0) );
fim FAN_N7057_1 ( .fault(fault), .net(N7057), .FEN(FEN[2731]), .op(N7057_t1) );
fim FAN_N7077_0 ( .fault(fault), .net(N7077), .FEN(FEN[2732]), .op(N7077_t0) );
fim FAN_N7077_1 ( .fault(fault), .net(N7077), .FEN(FEN[2733]), .op(N7077_t1) );
fim FAN_N7073_0 ( .fault(fault), .net(N7073), .FEN(FEN[2734]), .op(N7073_t0) );
fim FAN_N7073_1 ( .fault(fault), .net(N7073), .FEN(FEN[2735]), .op(N7073_t1) );
fim FAN_N7073_2 ( .fault(fault), .net(N7073), .FEN(FEN[2736]), .op(N7073_t2) );
fim FAN_N7068_0 ( .fault(fault), .net(N7068), .FEN(FEN[2737]), .op(N7068_t0) );
fim FAN_N7068_1 ( .fault(fault), .net(N7068), .FEN(FEN[2738]), .op(N7068_t1) );
fim FAN_N7068_2 ( .fault(fault), .net(N7068), .FEN(FEN[2739]), .op(N7068_t2) );
fim FAN_N7068_3 ( .fault(fault), .net(N7068), .FEN(FEN[2740]), .op(N7068_t3) );
fim FAN_N7095_0 ( .fault(fault), .net(N7095), .FEN(FEN[2741]), .op(N7095_t0) );
fim FAN_N7095_1 ( .fault(fault), .net(N7095), .FEN(FEN[2742]), .op(N7095_t1) );
fim FAN_N7091_0 ( .fault(fault), .net(N7091), .FEN(FEN[2743]), .op(N7091_t0) );
fim FAN_N7091_1 ( .fault(fault), .net(N7091), .FEN(FEN[2744]), .op(N7091_t1) );
fim FAN_N7091_2 ( .fault(fault), .net(N7091), .FEN(FEN[2745]), .op(N7091_t2) );
fim FAN_N7086_0 ( .fault(fault), .net(N7086), .FEN(FEN[2746]), .op(N7086_t0) );
fim FAN_N7086_1 ( .fault(fault), .net(N7086), .FEN(FEN[2747]), .op(N7086_t1) );
fim FAN_N7086_2 ( .fault(fault), .net(N7086), .FEN(FEN[2748]), .op(N7086_t2) );
fim FAN_N7086_3 ( .fault(fault), .net(N7086), .FEN(FEN[2749]), .op(N7086_t3) );
fim FAN_N7080_0 ( .fault(fault), .net(N7080), .FEN(FEN[2750]), .op(N7080_t0) );
fim FAN_N7080_1 ( .fault(fault), .net(N7080), .FEN(FEN[2751]), .op(N7080_t1) );
fim FAN_N7080_2 ( .fault(fault), .net(N7080), .FEN(FEN[2752]), .op(N7080_t2) );
fim FAN_N7080_3 ( .fault(fault), .net(N7080), .FEN(FEN[2753]), .op(N7080_t3) );
fim FAN_N7080_4 ( .fault(fault), .net(N7080), .FEN(FEN[2754]), .op(N7080_t4) );
fim FAN_N7100_0 ( .fault(fault), .net(N7100), .FEN(FEN[2755]), .op(N7100_t0) );
fim FAN_N7100_1 ( .fault(fault), .net(N7100), .FEN(FEN[2756]), .op(N7100_t1) );
fim FAN_N7114_0 ( .fault(fault), .net(N7114), .FEN(FEN[2757]), .op(N7114_t0) );
fim FAN_N7114_1 ( .fault(fault), .net(N7114), .FEN(FEN[2758]), .op(N7114_t1) );
fim FAN_N7114_2 ( .fault(fault), .net(N7114), .FEN(FEN[2759]), .op(N7114_t2) );
fim FAN_N7114_3 ( .fault(fault), .net(N7114), .FEN(FEN[2760]), .op(N7114_t3) );
fim FAN_N7114_4 ( .fault(fault), .net(N7114), .FEN(FEN[2761]), .op(N7114_t4) );
fim FAN_N7114_5 ( .fault(fault), .net(N7114), .FEN(FEN[2762]), .op(N7114_t5) );
fim FAN_N7114_6 ( .fault(fault), .net(N7114), .FEN(FEN[2763]), .op(N7114_t6) );
fim FAN_N7114_7 ( .fault(fault), .net(N7114), .FEN(FEN[2764]), .op(N7114_t7) );
fim FAN_N7114_8 ( .fault(fault), .net(N7114), .FEN(FEN[2765]), .op(N7114_t8) );
fim FAN_N7114_9 ( .fault(fault), .net(N7114), .FEN(FEN[2766]), .op(N7114_t9) );
fim FAN_N7125_0 ( .fault(fault), .net(N7125), .FEN(FEN[2767]), .op(N7125_t0) );
fim FAN_N7125_1 ( .fault(fault), .net(N7125), .FEN(FEN[2768]), .op(N7125_t1) );
fim FAN_N7125_2 ( .fault(fault), .net(N7125), .FEN(FEN[2769]), .op(N7125_t2) );
fim FAN_N7125_3 ( .fault(fault), .net(N7125), .FEN(FEN[2770]), .op(N7125_t3) );
fim FAN_N7125_4 ( .fault(fault), .net(N7125), .FEN(FEN[2771]), .op(N7125_t4) );
fim FAN_N7125_5 ( .fault(fault), .net(N7125), .FEN(FEN[2772]), .op(N7125_t5) );
fim FAN_N7125_6 ( .fault(fault), .net(N7125), .FEN(FEN[2773]), .op(N7125_t6) );
fim FAN_N7125_7 ( .fault(fault), .net(N7125), .FEN(FEN[2774]), .op(N7125_t7) );
fim FAN_N7125_8 ( .fault(fault), .net(N7125), .FEN(FEN[2775]), .op(N7125_t8) );
fim FAN_N7125_9 ( .fault(fault), .net(N7125), .FEN(FEN[2776]), .op(N7125_t9) );
fim FAN_N7107_0 ( .fault(fault), .net(N7107), .FEN(FEN[2777]), .op(N7107_t0) );
fim FAN_N7107_1 ( .fault(fault), .net(N7107), .FEN(FEN[2778]), .op(N7107_t1) );
fim FAN_N7107_2 ( .fault(fault), .net(N7107), .FEN(FEN[2779]), .op(N7107_t2) );
fim FAN_N7107_3 ( .fault(fault), .net(N7107), .FEN(FEN[2780]), .op(N7107_t3) );
fim FAN_N7107_4 ( .fault(fault), .net(N7107), .FEN(FEN[2781]), .op(N7107_t4) );
fim FAN_N7107_5 ( .fault(fault), .net(N7107), .FEN(FEN[2782]), .op(N7107_t5) );
fim FAN_N4657_0 ( .fault(fault), .net(N4657), .FEN(FEN[2783]), .op(N4657_t0) );
fim FAN_N4657_1 ( .fault(fault), .net(N4657), .FEN(FEN[2784]), .op(N4657_t1) );
fim FAN_N4657_2 ( .fault(fault), .net(N4657), .FEN(FEN[2785]), .op(N4657_t2) );
fim FAN_N4661_0 ( .fault(fault), .net(N4661), .FEN(FEN[2786]), .op(N4661_t0) );
fim FAN_N4661_1 ( .fault(fault), .net(N4661), .FEN(FEN[2787]), .op(N4661_t1) );
fim FAN_N4661_2 ( .fault(fault), .net(N4661), .FEN(FEN[2788]), .op(N4661_t2) );
fim FAN_N4661_3 ( .fault(fault), .net(N4661), .FEN(FEN[2789]), .op(N4661_t3) );
fim FAN_N4661_4 ( .fault(fault), .net(N4661), .FEN(FEN[2790]), .op(N4661_t4) );
fim FAN_N7149_0 ( .fault(fault), .net(N7149), .FEN(FEN[2791]), .op(N7149_t0) );
fim FAN_N7149_1 ( .fault(fault), .net(N7149), .FEN(FEN[2792]), .op(N7149_t1) );
fim FAN_N7149_2 ( .fault(fault), .net(N7149), .FEN(FEN[2793]), .op(N7149_t2) );
fim FAN_N7149_3 ( .fault(fault), .net(N7149), .FEN(FEN[2794]), .op(N7149_t3) );
fim FAN_N7149_4 ( .fault(fault), .net(N7149), .FEN(FEN[2795]), .op(N7149_t4) );
fim FAN_N7149_5 ( .fault(fault), .net(N7149), .FEN(FEN[2796]), .op(N7149_t5) );
fim FAN_N7149_6 ( .fault(fault), .net(N7149), .FEN(FEN[2797]), .op(N7149_t6) );
fim FAN_N7149_7 ( .fault(fault), .net(N7149), .FEN(FEN[2798]), .op(N7149_t7) );
fim FAN_N7149_8 ( .fault(fault), .net(N7149), .FEN(FEN[2799]), .op(N7149_t8) );
fim FAN_N7180_0 ( .fault(fault), .net(N7180), .FEN(FEN[2800]), .op(N7180_t0) );
fim FAN_N7180_1 ( .fault(fault), .net(N7180), .FEN(FEN[2801]), .op(N7180_t1) );
fim FAN_N7180_2 ( .fault(fault), .net(N7180), .FEN(FEN[2802]), .op(N7180_t2) );
fim FAN_N7180_3 ( .fault(fault), .net(N7180), .FEN(FEN[2803]), .op(N7180_t3) );
fim FAN_N7180_4 ( .fault(fault), .net(N7180), .FEN(FEN[2804]), .op(N7180_t4) );
fim FAN_N7180_5 ( .fault(fault), .net(N7180), .FEN(FEN[2805]), .op(N7180_t5) );
fim FAN_N7159_0 ( .fault(fault), .net(N7159), .FEN(FEN[2806]), .op(N7159_t0) );
fim FAN_N7159_1 ( .fault(fault), .net(N7159), .FEN(FEN[2807]), .op(N7159_t1) );
fim FAN_N7159_2 ( .fault(fault), .net(N7159), .FEN(FEN[2808]), .op(N7159_t2) );
fim FAN_N7159_3 ( .fault(fault), .net(N7159), .FEN(FEN[2809]), .op(N7159_t3) );
fim FAN_N7159_4 ( .fault(fault), .net(N7159), .FEN(FEN[2810]), .op(N7159_t4) );
fim FAN_N7159_5 ( .fault(fault), .net(N7159), .FEN(FEN[2811]), .op(N7159_t5) );
fim FAN_N7159_6 ( .fault(fault), .net(N7159), .FEN(FEN[2812]), .op(N7159_t6) );
fim FAN_N7159_7 ( .fault(fault), .net(N7159), .FEN(FEN[2813]), .op(N7159_t7) );
fim FAN_N7159_8 ( .fault(fault), .net(N7159), .FEN(FEN[2814]), .op(N7159_t8) );
fim FAN_N7159_9 ( .fault(fault), .net(N7159), .FEN(FEN[2815]), .op(N7159_t9) );
fim FAN_N7142_0 ( .fault(fault), .net(N7142), .FEN(FEN[2816]), .op(N7142_t0) );
fim FAN_N7142_1 ( .fault(fault), .net(N7142), .FEN(FEN[2817]), .op(N7142_t1) );
fim FAN_N7142_2 ( .fault(fault), .net(N7142), .FEN(FEN[2818]), .op(N7142_t2) );
fim FAN_N7142_3 ( .fault(fault), .net(N7142), .FEN(FEN[2819]), .op(N7142_t3) );
fim FAN_N7142_4 ( .fault(fault), .net(N7142), .FEN(FEN[2820]), .op(N7142_t4) );
fim FAN_N7142_5 ( .fault(fault), .net(N7142), .FEN(FEN[2821]), .op(N7142_t5) );
fim FAN_N7170_0 ( .fault(fault), .net(N7170), .FEN(FEN[2822]), .op(N7170_t0) );
fim FAN_N7170_1 ( .fault(fault), .net(N7170), .FEN(FEN[2823]), .op(N7170_t1) );
fim FAN_N7170_2 ( .fault(fault), .net(N7170), .FEN(FEN[2824]), .op(N7170_t2) );
fim FAN_N7170_3 ( .fault(fault), .net(N7170), .FEN(FEN[2825]), .op(N7170_t3) );
fim FAN_N7170_4 ( .fault(fault), .net(N7170), .FEN(FEN[2826]), .op(N7170_t4) );
fim FAN_N7170_5 ( .fault(fault), .net(N7170), .FEN(FEN[2827]), .op(N7170_t5) );
fim FAN_N7170_6 ( .fault(fault), .net(N7170), .FEN(FEN[2828]), .op(N7170_t6) );
fim FAN_N7170_7 ( .fault(fault), .net(N7170), .FEN(FEN[2829]), .op(N7170_t7) );
fim FAN_N7170_8 ( .fault(fault), .net(N7170), .FEN(FEN[2830]), .op(N7170_t8) );
fim FAN_N4675_0 ( .fault(fault), .net(N4675), .FEN(FEN[2831]), .op(N4675_t0) );
fim FAN_N4675_1 ( .fault(fault), .net(N4675), .FEN(FEN[2832]), .op(N4675_t1) );
fim FAN_N4678_0 ( .fault(fault), .net(N4678), .FEN(FEN[2833]), .op(N4678_t0) );
fim FAN_N4678_1 ( .fault(fault), .net(N4678), .FEN(FEN[2834]), .op(N4678_t1) );
fim FAN_N4678_2 ( .fault(fault), .net(N4678), .FEN(FEN[2835]), .op(N4678_t2) );
fim FAN_N4682_0 ( .fault(fault), .net(N4682), .FEN(FEN[2836]), .op(N4682_t0) );
fim FAN_N4682_1 ( .fault(fault), .net(N4682), .FEN(FEN[2837]), .op(N4682_t1) );
fim FAN_N4682_2 ( .fault(fault), .net(N4682), .FEN(FEN[2838]), .op(N4682_t2) );
fim FAN_N4682_3 ( .fault(fault), .net(N4682), .FEN(FEN[2839]), .op(N4682_t3) );
fim FAN_N4687_0 ( .fault(fault), .net(N4687), .FEN(FEN[2840]), .op(N4687_t0) );
fim FAN_N4687_1 ( .fault(fault), .net(N4687), .FEN(FEN[2841]), .op(N4687_t1) );
fim FAN_N4687_2 ( .fault(fault), .net(N4687), .FEN(FEN[2842]), .op(N4687_t2) );
fim FAN_N4687_3 ( .fault(fault), .net(N4687), .FEN(FEN[2843]), .op(N4687_t3) );
fim FAN_N4687_4 ( .fault(fault), .net(N4687), .FEN(FEN[2844]), .op(N4687_t4) );
fim FAN_N7194_0 ( .fault(fault), .net(N7194), .FEN(FEN[2845]), .op(N7194_t0) );
fim FAN_N7194_1 ( .fault(fault), .net(N7194), .FEN(FEN[2846]), .op(N7194_t1) );
fim FAN_N7194_2 ( .fault(fault), .net(N7194), .FEN(FEN[2847]), .op(N7194_t2) );
fim FAN_N7198_0 ( .fault(fault), .net(N7198), .FEN(FEN[2848]), .op(N7198_t0) );
fim FAN_N7198_1 ( .fault(fault), .net(N7198), .FEN(FEN[2849]), .op(N7198_t1) );
fim FAN_N7198_2 ( .fault(fault), .net(N7198), .FEN(FEN[2850]), .op(N7198_t2) );
fim FAN_N7205_0 ( .fault(fault), .net(N7205), .FEN(FEN[2851]), .op(N7205_t0) );
fim FAN_N7205_1 ( .fault(fault), .net(N7205), .FEN(FEN[2852]), .op(N7205_t1) );
fim FAN_N7205_2 ( .fault(fault), .net(N7205), .FEN(FEN[2853]), .op(N7205_t2) );
fim FAN_N7209_0 ( .fault(fault), .net(N7209), .FEN(FEN[2854]), .op(N7209_t0) );
fim FAN_N7209_1 ( .fault(fault), .net(N7209), .FEN(FEN[2855]), .op(N7209_t1) );
fim FAN_N7209_2 ( .fault(fault), .net(N7209), .FEN(FEN[2856]), .op(N7209_t2) );
fim FAN_N7216_0 ( .fault(fault), .net(N7216), .FEN(FEN[2857]), .op(N7216_t0) );
fim FAN_N7216_1 ( .fault(fault), .net(N7216), .FEN(FEN[2858]), .op(N7216_t1) );
fim FAN_N7219_0 ( .fault(fault), .net(N7219), .FEN(FEN[2859]), .op(N7219_t0) );
fim FAN_N7219_1 ( .fault(fault), .net(N7219), .FEN(FEN[2860]), .op(N7219_t1) );
fim FAN_N7202_0 ( .fault(fault), .net(N7202), .FEN(FEN[2861]), .op(N7202_t0) );
fim FAN_N7202_1 ( .fault(fault), .net(N7202), .FEN(FEN[2862]), .op(N7202_t1) );
fim FAN_N7213_0 ( .fault(fault), .net(N7213), .FEN(FEN[2863]), .op(N7213_t0) );
fim FAN_N7213_1 ( .fault(fault), .net(N7213), .FEN(FEN[2864]), .op(N7213_t1) );
fim FAN_N7191_0 ( .fault(fault), .net(N7191), .FEN(FEN[2865]), .op(N7191_t0) );
fim FAN_N7191_1 ( .fault(fault), .net(N7191), .FEN(FEN[2866]), .op(N7191_t1) );
fim FAN_N7188_0 ( .fault(fault), .net(N7188), .FEN(FEN[2867]), .op(N7188_t0) );
fim FAN_N7188_1 ( .fault(fault), .net(N7188), .FEN(FEN[2868]), .op(N7188_t1) );
fim FAN_N7301_0 ( .fault(fault), .net(N7301), .FEN(FEN[2869]), .op(N7301_t0) );
fim FAN_N7301_1 ( .fault(fault), .net(N7301), .FEN(FEN[2870]), .op(N7301_t1) );
fim FAN_N7301_2 ( .fault(fault), .net(N7301), .FEN(FEN[2871]), .op(N7301_t2) );
fim FAN_N7301_3 ( .fault(fault), .net(N7301), .FEN(FEN[2872]), .op(N7301_t3) );
fim FAN_N7301_4 ( .fault(fault), .net(N7301), .FEN(FEN[2873]), .op(N7301_t4) );
fim FAN_N7240_0 ( .fault(fault), .net(N7240), .FEN(FEN[2874]), .op(N7240_t0) );
fim FAN_N7240_1 ( .fault(fault), .net(N7240), .FEN(FEN[2875]), .op(N7240_t1) );
fim FAN_N7240_2 ( .fault(fault), .net(N7240), .FEN(FEN[2876]), .op(N7240_t2) );
fim FAN_N7240_3 ( .fault(fault), .net(N7240), .FEN(FEN[2877]), .op(N7240_t3) );
fim FAN_N7240_4 ( .fault(fault), .net(N7240), .FEN(FEN[2878]), .op(N7240_t4) );
fim FAN_N7240_5 ( .fault(fault), .net(N7240), .FEN(FEN[2879]), .op(N7240_t5) );
fim FAN_N7240_6 ( .fault(fault), .net(N7240), .FEN(FEN[2880]), .op(N7240_t6) );
fim FAN_N7240_7 ( .fault(fault), .net(N7240), .FEN(FEN[2881]), .op(N7240_t7) );
fim FAN_N7240_8 ( .fault(fault), .net(N7240), .FEN(FEN[2882]), .op(N7240_t8) );
fim FAN_N7229_0 ( .fault(fault), .net(N7229), .FEN(FEN[2883]), .op(N7229_t0) );
fim FAN_N7229_1 ( .fault(fault), .net(N7229), .FEN(FEN[2884]), .op(N7229_t1) );
fim FAN_N7229_2 ( .fault(fault), .net(N7229), .FEN(FEN[2885]), .op(N7229_t2) );
fim FAN_N7229_3 ( .fault(fault), .net(N7229), .FEN(FEN[2886]), .op(N7229_t3) );
fim FAN_N7229_4 ( .fault(fault), .net(N7229), .FEN(FEN[2887]), .op(N7229_t4) );
fim FAN_N7229_5 ( .fault(fault), .net(N7229), .FEN(FEN[2888]), .op(N7229_t5) );
fim FAN_N7229_6 ( .fault(fault), .net(N7229), .FEN(FEN[2889]), .op(N7229_t6) );
fim FAN_N7229_7 ( .fault(fault), .net(N7229), .FEN(FEN[2890]), .op(N7229_t7) );
fim FAN_N7229_8 ( .fault(fault), .net(N7229), .FEN(FEN[2891]), .op(N7229_t8) );
fim FAN_N7229_9 ( .fault(fault), .net(N7229), .FEN(FEN[2892]), .op(N7229_t9) );
fim FAN_N7222_0 ( .fault(fault), .net(N7222), .FEN(FEN[2893]), .op(N7222_t0) );
fim FAN_N7222_1 ( .fault(fault), .net(N7222), .FEN(FEN[2894]), .op(N7222_t1) );
fim FAN_N7222_2 ( .fault(fault), .net(N7222), .FEN(FEN[2895]), .op(N7222_t2) );
fim FAN_N7222_3 ( .fault(fault), .net(N7222), .FEN(FEN[2896]), .op(N7222_t3) );
fim FAN_N7222_4 ( .fault(fault), .net(N7222), .FEN(FEN[2897]), .op(N7222_t4) );
fim FAN_N7222_5 ( .fault(fault), .net(N7222), .FEN(FEN[2898]), .op(N7222_t5) );
fim FAN_N4702_0 ( .fault(fault), .net(N4702), .FEN(FEN[2899]), .op(N4702_t0) );
fim FAN_N4702_1 ( .fault(fault), .net(N4702), .FEN(FEN[2900]), .op(N4702_t1) );
fim FAN_N4702_2 ( .fault(fault), .net(N4702), .FEN(FEN[2901]), .op(N4702_t2) );
fim FAN_N4706_0 ( .fault(fault), .net(N4706), .FEN(FEN[2902]), .op(N4706_t0) );
fim FAN_N4706_1 ( .fault(fault), .net(N4706), .FEN(FEN[2903]), .op(N4706_t1) );
fim FAN_N4706_2 ( .fault(fault), .net(N4706), .FEN(FEN[2904]), .op(N4706_t2) );
fim FAN_N4706_3 ( .fault(fault), .net(N4706), .FEN(FEN[2905]), .op(N4706_t3) );
fim FAN_N7307_0 ( .fault(fault), .net(N7307), .FEN(FEN[2906]), .op(N7307_t0) );
fim FAN_N7307_1 ( .fault(fault), .net(N7307), .FEN(FEN[2907]), .op(N7307_t1) );
fim FAN_N7307_2 ( .fault(fault), .net(N7307), .FEN(FEN[2908]), .op(N7307_t2) );
fim FAN_N7307_3 ( .fault(fault), .net(N7307), .FEN(FEN[2909]), .op(N7307_t3) );
fim FAN_N7307_4 ( .fault(fault), .net(N7307), .FEN(FEN[2910]), .op(N7307_t4) );
fim FAN_N7307_5 ( .fault(fault), .net(N7307), .FEN(FEN[2911]), .op(N7307_t5) );
fim FAN_N7288_0 ( .fault(fault), .net(N7288), .FEN(FEN[2912]), .op(N7288_t0) );
fim FAN_N7288_1 ( .fault(fault), .net(N7288), .FEN(FEN[2913]), .op(N7288_t1) );
fim FAN_N7288_2 ( .fault(fault), .net(N7288), .FEN(FEN[2914]), .op(N7288_t2) );
fim FAN_N7288_3 ( .fault(fault), .net(N7288), .FEN(FEN[2915]), .op(N7288_t3) );
fim FAN_N7288_4 ( .fault(fault), .net(N7288), .FEN(FEN[2916]), .op(N7288_t4) );
fim FAN_N7288_5 ( .fault(fault), .net(N7288), .FEN(FEN[2917]), .op(N7288_t5) );
fim FAN_N7288_6 ( .fault(fault), .net(N7288), .FEN(FEN[2918]), .op(N7288_t6) );
fim FAN_N7288_7 ( .fault(fault), .net(N7288), .FEN(FEN[2919]), .op(N7288_t7) );
fim FAN_N7288_8 ( .fault(fault), .net(N7288), .FEN(FEN[2920]), .op(N7288_t8) );
fim FAN_N7288_9 ( .fault(fault), .net(N7288), .FEN(FEN[2921]), .op(N7288_t9) );
fim FAN_N7288_10 ( .fault(fault), .net(N7288), .FEN(FEN[2922]), .op(N7288_t10) );
fim FAN_N7288_11 ( .fault(fault), .net(N7288), .FEN(FEN[2923]), .op(N7288_t11) );
fim FAN_N7272_0 ( .fault(fault), .net(N7272), .FEN(FEN[2924]), .op(N7272_t0) );
fim FAN_N7272_1 ( .fault(fault), .net(N7272), .FEN(FEN[2925]), .op(N7272_t1) );
fim FAN_N7272_2 ( .fault(fault), .net(N7272), .FEN(FEN[2926]), .op(N7272_t2) );
fim FAN_N7272_3 ( .fault(fault), .net(N7272), .FEN(FEN[2927]), .op(N7272_t3) );
fim FAN_N7272_4 ( .fault(fault), .net(N7272), .FEN(FEN[2928]), .op(N7272_t4) );
fim FAN_N7272_5 ( .fault(fault), .net(N7272), .FEN(FEN[2929]), .op(N7272_t5) );
fim FAN_N7272_6 ( .fault(fault), .net(N7272), .FEN(FEN[2930]), .op(N7272_t6) );
fim FAN_N7272_7 ( .fault(fault), .net(N7272), .FEN(FEN[2931]), .op(N7272_t7) );
fim FAN_N7272_8 ( .fault(fault), .net(N7272), .FEN(FEN[2932]), .op(N7272_t8) );
fim FAN_N7272_9 ( .fault(fault), .net(N7272), .FEN(FEN[2933]), .op(N7272_t9) );
fim FAN_N7272_10 ( .fault(fault), .net(N7272), .FEN(FEN[2934]), .op(N7272_t10) );
fim FAN_N7272_11 ( .fault(fault), .net(N7272), .FEN(FEN[2935]), .op(N7272_t11) );
fim FAN_N7272_12 ( .fault(fault), .net(N7272), .FEN(FEN[2936]), .op(N7272_t12) );
fim FAN_N7272_13 ( .fault(fault), .net(N7272), .FEN(FEN[2937]), .op(N7272_t13) );
fim FAN_N7272_14 ( .fault(fault), .net(N7272), .FEN(FEN[2938]), .op(N7272_t14) );
fim FAN_N7258_0 ( .fault(fault), .net(N7258), .FEN(FEN[2939]), .op(N7258_t0) );
fim FAN_N7258_1 ( .fault(fault), .net(N7258), .FEN(FEN[2940]), .op(N7258_t1) );
fim FAN_N7258_2 ( .fault(fault), .net(N7258), .FEN(FEN[2941]), .op(N7258_t2) );
fim FAN_N7258_3 ( .fault(fault), .net(N7258), .FEN(FEN[2942]), .op(N7258_t3) );
fim FAN_N7258_4 ( .fault(fault), .net(N7258), .FEN(FEN[2943]), .op(N7258_t4) );
fim FAN_N7258_5 ( .fault(fault), .net(N7258), .FEN(FEN[2944]), .op(N7258_t5) );
fim FAN_N7258_6 ( .fault(fault), .net(N7258), .FEN(FEN[2945]), .op(N7258_t6) );
fim FAN_N7258_7 ( .fault(fault), .net(N7258), .FEN(FEN[2946]), .op(N7258_t7) );
fim FAN_N7258_8 ( .fault(fault), .net(N7258), .FEN(FEN[2947]), .op(N7258_t8) );
fim FAN_N7258_9 ( .fault(fault), .net(N7258), .FEN(FEN[2948]), .op(N7258_t9) );
fim FAN_N7258_10 ( .fault(fault), .net(N7258), .FEN(FEN[2949]), .op(N7258_t10) );
fim FAN_N7258_11 ( .fault(fault), .net(N7258), .FEN(FEN[2950]), .op(N7258_t11) );
fim FAN_N7258_12 ( .fault(fault), .net(N7258), .FEN(FEN[2951]), .op(N7258_t12) );
fim FAN_N7250_0 ( .fault(fault), .net(N7250), .FEN(FEN[2952]), .op(N7250_t0) );
fim FAN_N7250_1 ( .fault(fault), .net(N7250), .FEN(FEN[2953]), .op(N7250_t1) );
fim FAN_N7250_2 ( .fault(fault), .net(N7250), .FEN(FEN[2954]), .op(N7250_t2) );
fim FAN_N7250_3 ( .fault(fault), .net(N7250), .FEN(FEN[2955]), .op(N7250_t3) );
fim FAN_N7250_4 ( .fault(fault), .net(N7250), .FEN(FEN[2956]), .op(N7250_t4) );
fim FAN_N7250_5 ( .fault(fault), .net(N7250), .FEN(FEN[2957]), .op(N7250_t5) );
fim FAN_N7250_6 ( .fault(fault), .net(N7250), .FEN(FEN[2958]), .op(N7250_t6) );
fim FAN_N4718_0 ( .fault(fault), .net(N4718), .FEN(FEN[2959]), .op(N4718_t0) );
fim FAN_N4718_1 ( .fault(fault), .net(N4718), .FEN(FEN[2960]), .op(N4718_t1) );
fim FAN_N4718_2 ( .fault(fault), .net(N4718), .FEN(FEN[2961]), .op(N4718_t2) );
fim FAN_N4722_0 ( .fault(fault), .net(N4722), .FEN(FEN[2962]), .op(N4722_t0) );
fim FAN_N4722_1 ( .fault(fault), .net(N4722), .FEN(FEN[2963]), .op(N4722_t1) );
fim FAN_N4722_2 ( .fault(fault), .net(N4722), .FEN(FEN[2964]), .op(N4722_t2) );
fim FAN_N4722_3 ( .fault(fault), .net(N4722), .FEN(FEN[2965]), .op(N4722_t3) );
fim FAN_N4722_4 ( .fault(fault), .net(N4722), .FEN(FEN[2966]), .op(N4722_t4) );
fim FAN_N4728_0 ( .fault(fault), .net(N4728), .FEN(FEN[2967]), .op(N4728_t0) );
fim FAN_N4728_1 ( .fault(fault), .net(N4728), .FEN(FEN[2968]), .op(N4728_t1) );
fim FAN_N4728_2 ( .fault(fault), .net(N4728), .FEN(FEN[2969]), .op(N4728_t2) );
fim FAN_N4728_3 ( .fault(fault), .net(N4728), .FEN(FEN[2970]), .op(N4728_t3) );
fim FAN_N4728_4 ( .fault(fault), .net(N4728), .FEN(FEN[2971]), .op(N4728_t4) );
fim FAN_N4728_5 ( .fault(fault), .net(N4728), .FEN(FEN[2972]), .op(N4728_t5) );
fim FAN_N7314_0 ( .fault(fault), .net(N7314), .FEN(FEN[2973]), .op(N7314_t0) );
fim FAN_N7314_1 ( .fault(fault), .net(N7314), .FEN(FEN[2974]), .op(N7314_t1) );
fim FAN_N7314_2 ( .fault(fault), .net(N7314), .FEN(FEN[2975]), .op(N7314_t2) );
fim FAN_N7318_0 ( .fault(fault), .net(N7318), .FEN(FEN[2976]), .op(N7318_t0) );
fim FAN_N7318_1 ( .fault(fault), .net(N7318), .FEN(FEN[2977]), .op(N7318_t1) );
fim FAN_N7318_2 ( .fault(fault), .net(N7318), .FEN(FEN[2978]), .op(N7318_t2) );
fim FAN_N7322_0 ( .fault(fault), .net(N7322), .FEN(FEN[2979]), .op(N7322_t0) );
fim FAN_N7322_1 ( .fault(fault), .net(N7322), .FEN(FEN[2980]), .op(N7322_t1) );
fim FAN_N7331_0 ( .fault(fault), .net(N7331), .FEN(FEN[2981]), .op(N7331_t0) );
fim FAN_N7331_1 ( .fault(fault), .net(N7331), .FEN(FEN[2982]), .op(N7331_t1) );
fim FAN_N7340_0 ( .fault(fault), .net(N7340), .FEN(FEN[2983]), .op(N7340_t0) );
fim FAN_N7340_1 ( .fault(fault), .net(N7340), .FEN(FEN[2984]), .op(N7340_t1) );
fim FAN_N7343_0 ( .fault(fault), .net(N7343), .FEN(FEN[2985]), .op(N7343_t0) );
fim FAN_N7343_1 ( .fault(fault), .net(N7343), .FEN(FEN[2986]), .op(N7343_t1) );
fim FAN_N7337_0 ( .fault(fault), .net(N7337), .FEN(FEN[2987]), .op(N7337_t0) );
fim FAN_N7337_1 ( .fault(fault), .net(N7337), .FEN(FEN[2988]), .op(N7337_t1) );
fim FAN_N7334_0 ( .fault(fault), .net(N7334), .FEN(FEN[2989]), .op(N7334_t0) );
fim FAN_N7334_1 ( .fault(fault), .net(N7334), .FEN(FEN[2990]), .op(N7334_t1) );
fim FAN_N7355_0 ( .fault(fault), .net(N7355), .FEN(FEN[2991]), .op(N7355_t0) );
fim FAN_N7355_1 ( .fault(fault), .net(N7355), .FEN(FEN[2992]), .op(N7355_t1) );
fim FAN_N7351_0 ( .fault(fault), .net(N7351), .FEN(FEN[2993]), .op(N7351_t0) );
fim FAN_N7351_1 ( .fault(fault), .net(N7351), .FEN(FEN[2994]), .op(N7351_t1) );
fim FAN_N7351_2 ( .fault(fault), .net(N7351), .FEN(FEN[2995]), .op(N7351_t2) );
fim FAN_N7346_0 ( .fault(fault), .net(N7346), .FEN(FEN[2996]), .op(N7346_t0) );
fim FAN_N7346_1 ( .fault(fault), .net(N7346), .FEN(FEN[2997]), .op(N7346_t1) );
fim FAN_N7346_2 ( .fault(fault), .net(N7346), .FEN(FEN[2998]), .op(N7346_t2) );
fim FAN_N7346_3 ( .fault(fault), .net(N7346), .FEN(FEN[2999]), .op(N7346_t3) );
fim FAN_N7373_0 ( .fault(fault), .net(N7373), .FEN(FEN[3000]), .op(N7373_t0) );
fim FAN_N7373_1 ( .fault(fault), .net(N7373), .FEN(FEN[3001]), .op(N7373_t1) );
fim FAN_N7369_0 ( .fault(fault), .net(N7369), .FEN(FEN[3002]), .op(N7369_t0) );
fim FAN_N7369_1 ( .fault(fault), .net(N7369), .FEN(FEN[3003]), .op(N7369_t1) );
fim FAN_N7369_2 ( .fault(fault), .net(N7369), .FEN(FEN[3004]), .op(N7369_t2) );
fim FAN_N7364_0 ( .fault(fault), .net(N7364), .FEN(FEN[3005]), .op(N7364_t0) );
fim FAN_N7364_1 ( .fault(fault), .net(N7364), .FEN(FEN[3006]), .op(N7364_t1) );
fim FAN_N7364_2 ( .fault(fault), .net(N7364), .FEN(FEN[3007]), .op(N7364_t2) );
fim FAN_N7364_3 ( .fault(fault), .net(N7364), .FEN(FEN[3008]), .op(N7364_t3) );
fim FAN_N7358_0 ( .fault(fault), .net(N7358), .FEN(FEN[3009]), .op(N7358_t0) );
fim FAN_N7358_1 ( .fault(fault), .net(N7358), .FEN(FEN[3010]), .op(N7358_t1) );
fim FAN_N7358_2 ( .fault(fault), .net(N7358), .FEN(FEN[3011]), .op(N7358_t2) );
fim FAN_N7358_3 ( .fault(fault), .net(N7358), .FEN(FEN[3012]), .op(N7358_t3) );
fim FAN_N7358_4 ( .fault(fault), .net(N7358), .FEN(FEN[3013]), .op(N7358_t4) );
fim FAN_N7387_0 ( .fault(fault), .net(N7387), .FEN(FEN[3014]), .op(N7387_t0) );
fim FAN_N7387_1 ( .fault(fault), .net(N7387), .FEN(FEN[3015]), .op(N7387_t1) );
fim FAN_N7387_2 ( .fault(fault), .net(N7387), .FEN(FEN[3016]), .op(N7387_t2) );
fim FAN_N7394_0 ( .fault(fault), .net(N7394), .FEN(FEN[3017]), .op(N7394_t0) );
fim FAN_N7394_1 ( .fault(fault), .net(N7394), .FEN(FEN[3018]), .op(N7394_t1) );
fim FAN_N7394_2 ( .fault(fault), .net(N7394), .FEN(FEN[3019]), .op(N7394_t2) );
fim FAN_N7398_0 ( .fault(fault), .net(N7398), .FEN(FEN[3020]), .op(N7398_t0) );
fim FAN_N7398_1 ( .fault(fault), .net(N7398), .FEN(FEN[3021]), .op(N7398_t1) );
fim FAN_N7398_2 ( .fault(fault), .net(N7398), .FEN(FEN[3022]), .op(N7398_t2) );
fim FAN_N7405_0 ( .fault(fault), .net(N7405), .FEN(FEN[3023]), .op(N7405_t0) );
fim FAN_N7405_1 ( .fault(fault), .net(N7405), .FEN(FEN[3024]), .op(N7405_t1) );
fim FAN_N7408_0 ( .fault(fault), .net(N7408), .FEN(FEN[3025]), .op(N7408_t0) );
fim FAN_N7408_1 ( .fault(fault), .net(N7408), .FEN(FEN[3026]), .op(N7408_t1) );
fim FAN_N7391_0 ( .fault(fault), .net(N7391), .FEN(FEN[3027]), .op(N7391_t0) );
fim FAN_N7391_1 ( .fault(fault), .net(N7391), .FEN(FEN[3028]), .op(N7391_t1) );
fim FAN_N7402_0 ( .fault(fault), .net(N7402), .FEN(FEN[3029]), .op(N7402_t0) );
fim FAN_N7402_1 ( .fault(fault), .net(N7402), .FEN(FEN[3030]), .op(N7402_t1) );
fim FAN_N7381_0 ( .fault(fault), .net(N7381), .FEN(FEN[3031]), .op(N7381_t0) );
fim FAN_N7381_1 ( .fault(fault), .net(N7381), .FEN(FEN[3032]), .op(N7381_t1) );
fim FAN_N7378_0 ( .fault(fault), .net(N7378), .FEN(FEN[3033]), .op(N7378_t0) );
fim FAN_N7378_1 ( .fault(fault), .net(N7378), .FEN(FEN[3034]), .op(N7378_t1) );
fim FAN_N7441_0 ( .fault(fault), .net(N7441), .FEN(FEN[3035]), .op(N7441_t0) );
fim FAN_N7441_1 ( .fault(fault), .net(N7441), .FEN(FEN[3036]), .op(N7441_t1) );
fim FAN_N7444_0 ( .fault(fault), .net(N7444), .FEN(FEN[3037]), .op(N7444_t0) );
fim FAN_N7444_1 ( .fault(fault), .net(N7444), .FEN(FEN[3038]), .op(N7444_t1) );
fim FAN_N7447_0 ( .fault(fault), .net(N7447), .FEN(FEN[3039]), .op(N7447_t0) );
fim FAN_N7447_1 ( .fault(fault), .net(N7447), .FEN(FEN[3040]), .op(N7447_t1) );
fim FAN_N7450_0 ( .fault(fault), .net(N7450), .FEN(FEN[3041]), .op(N7450_t0) );
fim FAN_N7450_1 ( .fault(fault), .net(N7450), .FEN(FEN[3042]), .op(N7450_t1) );
fim FAN_N7453_0 ( .fault(fault), .net(N7453), .FEN(FEN[3043]), .op(N7453_t0) );
fim FAN_N7453_1 ( .fault(fault), .net(N7453), .FEN(FEN[3044]), .op(N7453_t1) );
fim FAN_N7456_0 ( .fault(fault), .net(N7456), .FEN(FEN[3045]), .op(N7456_t0) );
fim FAN_N7456_1 ( .fault(fault), .net(N7456), .FEN(FEN[3046]), .op(N7456_t1) );
fim FAN_N7474_0 ( .fault(fault), .net(N7474), .FEN(FEN[3047]), .op(N7474_t0) );
fim FAN_N7474_1 ( .fault(fault), .net(N7474), .FEN(FEN[3048]), .op(N7474_t1) );
fim FAN_N7465_0 ( .fault(fault), .net(N7465), .FEN(FEN[3049]), .op(N7465_t0) );
fim FAN_N7465_1 ( .fault(fault), .net(N7465), .FEN(FEN[3050]), .op(N7465_t1) );
fim FAN_N7468_0 ( .fault(fault), .net(N7468), .FEN(FEN[3051]), .op(N7468_t0) );
fim FAN_N7468_1 ( .fault(fault), .net(N7468), .FEN(FEN[3052]), .op(N7468_t1) );
fim FAN_N7471_0 ( .fault(fault), .net(N7471), .FEN(FEN[3053]), .op(N7471_t0) );
fim FAN_N7471_1 ( .fault(fault), .net(N7471), .FEN(FEN[3054]), .op(N7471_t1) );
fim FAN_N7479_0 ( .fault(fault), .net(N7479), .FEN(FEN[3055]), .op(N7479_t0) );
fim FAN_N7479_1 ( .fault(fault), .net(N7479), .FEN(FEN[3056]), .op(N7479_t1) );
fim FAN_N7482_0 ( .fault(fault), .net(N7482), .FEN(FEN[3057]), .op(N7482_t0) );
fim FAN_N7482_1 ( .fault(fault), .net(N7482), .FEN(FEN[3058]), .op(N7482_t1) );
fim FAN_N7485_0 ( .fault(fault), .net(N7485), .FEN(FEN[3059]), .op(N7485_t0) );
fim FAN_N7485_1 ( .fault(fault), .net(N7485), .FEN(FEN[3060]), .op(N7485_t1) );
fim FAN_N7491_0 ( .fault(fault), .net(N7491), .FEN(FEN[3061]), .op(N7491_t0) );
fim FAN_N7491_1 ( .fault(fault), .net(N7491), .FEN(FEN[3062]), .op(N7491_t1) );
fim FAN_N7494_0 ( .fault(fault), .net(N7494), .FEN(FEN[3063]), .op(N7494_t0) );
fim FAN_N7494_1 ( .fault(fault), .net(N7494), .FEN(FEN[3064]), .op(N7494_t1) );
fim FAN_N7497_0 ( .fault(fault), .net(N7497), .FEN(FEN[3065]), .op(N7497_t0) );
fim FAN_N7497_1 ( .fault(fault), .net(N7497), .FEN(FEN[3066]), .op(N7497_t1) );
fim FAN_N7503_0 ( .fault(fault), .net(N7503), .FEN(FEN[3067]), .op(N7503_t0) );
fim FAN_N7503_1 ( .fault(fault), .net(N7503), .FEN(FEN[3068]), .op(N7503_t1) );
fim FAN_N7506_0 ( .fault(fault), .net(N7506), .FEN(FEN[3069]), .op(N7506_t0) );
fim FAN_N7506_1 ( .fault(fault), .net(N7506), .FEN(FEN[3070]), .op(N7506_t1) );
fim FAN_N7509_0 ( .fault(fault), .net(N7509), .FEN(FEN[3071]), .op(N7509_t0) );
fim FAN_N7509_1 ( .fault(fault), .net(N7509), .FEN(FEN[3072]), .op(N7509_t1) );
fim FAN_N7512_0 ( .fault(fault), .net(N7512), .FEN(FEN[3073]), .op(N7512_t0) );
fim FAN_N7512_1 ( .fault(fault), .net(N7512), .FEN(FEN[3074]), .op(N7512_t1) );
fim FAN_N7530_0 ( .fault(fault), .net(N7530), .FEN(FEN[3075]), .op(N7530_t0) );
fim FAN_N7530_1 ( .fault(fault), .net(N7530), .FEN(FEN[3076]), .op(N7530_t1) );
fim FAN_N7521_0 ( .fault(fault), .net(N7521), .FEN(FEN[3077]), .op(N7521_t0) );
fim FAN_N7521_1 ( .fault(fault), .net(N7521), .FEN(FEN[3078]), .op(N7521_t1) );
fim FAN_N7524_0 ( .fault(fault), .net(N7524), .FEN(FEN[3079]), .op(N7524_t0) );
fim FAN_N7524_1 ( .fault(fault), .net(N7524), .FEN(FEN[3080]), .op(N7524_t1) );
fim FAN_N7527_0 ( .fault(fault), .net(N7527), .FEN(FEN[3081]), .op(N7527_t0) );
fim FAN_N7527_1 ( .fault(fault), .net(N7527), .FEN(FEN[3082]), .op(N7527_t1) );
fim FAN_N7553_0 ( .fault(fault), .net(N7553), .FEN(FEN[3083]), .op(N7553_t0) );
fim FAN_N7553_1 ( .fault(fault), .net(N7553), .FEN(FEN[3084]), .op(N7553_t1) );
fim FAN_N7574_0 ( .fault(fault), .net(N7574), .FEN(FEN[3085]), .op(N7574_t0) );
fim FAN_N7574_1 ( .fault(fault), .net(N7574), .FEN(FEN[3086]), .op(N7574_t1) );
fim FAN_N7577_0 ( .fault(fault), .net(N7577), .FEN(FEN[3087]), .op(N7577_t0) );
fim FAN_N7577_1 ( .fault(fault), .net(N7577), .FEN(FEN[3088]), .op(N7577_t1) );
fim FAN_N7560_0 ( .fault(fault), .net(N7560), .FEN(FEN[3089]), .op(N7560_t0) );
fim FAN_N7560_1 ( .fault(fault), .net(N7560), .FEN(FEN[3090]), .op(N7560_t1) );
fim FAN_N7563_0 ( .fault(fault), .net(N7563), .FEN(FEN[3091]), .op(N7563_t0) );
fim FAN_N7563_1 ( .fault(fault), .net(N7563), .FEN(FEN[3092]), .op(N7563_t1) );
fim FAN_N7566_0 ( .fault(fault), .net(N7566), .FEN(FEN[3093]), .op(N7566_t0) );
fim FAN_N7566_1 ( .fault(fault), .net(N7566), .FEN(FEN[3094]), .op(N7566_t1) );
fim FAN_N7569_0 ( .fault(fault), .net(N7569), .FEN(FEN[3095]), .op(N7569_t0) );
fim FAN_N7569_1 ( .fault(fault), .net(N7569), .FEN(FEN[3096]), .op(N7569_t1) );
fim FAN_N7588_0 ( .fault(fault), .net(N7588), .FEN(FEN[3097]), .op(N7588_t0) );
fim FAN_N7588_1 ( .fault(fault), .net(N7588), .FEN(FEN[3098]), .op(N7588_t1) );
fim FAN_N7591_0 ( .fault(fault), .net(N7591), .FEN(FEN[3099]), .op(N7591_t0) );
fim FAN_N7591_1 ( .fault(fault), .net(N7591), .FEN(FEN[3100]), .op(N7591_t1) );
fim FAN_N7582_0 ( .fault(fault), .net(N7582), .FEN(FEN[3101]), .op(N7582_t0) );
fim FAN_N7582_1 ( .fault(fault), .net(N7582), .FEN(FEN[3102]), .op(N7582_t1) );
fim FAN_N7585_0 ( .fault(fault), .net(N7585), .FEN(FEN[3103]), .op(N7585_t0) );
fim FAN_N7585_1 ( .fault(fault), .net(N7585), .FEN(FEN[3104]), .op(N7585_t1) );
fim FAN_N7620_0 ( .fault(fault), .net(N7620), .FEN(FEN[3105]), .op(N7620_t0) );
fim FAN_N7620_1 ( .fault(fault), .net(N7620), .FEN(FEN[3106]), .op(N7620_t1) );
fim FAN_N7609_0 ( .fault(fault), .net(N7609), .FEN(FEN[3107]), .op(N7609_t0) );
fim FAN_N7609_1 ( .fault(fault), .net(N7609), .FEN(FEN[3108]), .op(N7609_t1) );
fim FAN_N7609_2 ( .fault(fault), .net(N7609), .FEN(FEN[3109]), .op(N7609_t2) );
fim FAN_N7655_0 ( .fault(fault), .net(N7655), .FEN(FEN[3110]), .op(N7655_t0) );
fim FAN_N7655_1 ( .fault(fault), .net(N7655), .FEN(FEN[3111]), .op(N7655_t1) );
fim FAN_N7655_2 ( .fault(fault), .net(N7655), .FEN(FEN[3112]), .op(N7655_t2) );
fim FAN_N7671_0 ( .fault(fault), .net(N7671), .FEN(FEN[3113]), .op(N7671_t0) );
fim FAN_N7671_1 ( .fault(fault), .net(N7671), .FEN(FEN[3114]), .op(N7671_t1) );
fim FAN_N8196_0 ( .fault(fault), .net(N8196), .FEN(FEN[3115]), .op(N8196_t0) );
fim FAN_N8196_1 ( .fault(fault), .net(N8196), .FEN(FEN[3116]), .op(N8196_t1) );
fim FAN_N8200_0 ( .fault(fault), .net(N8200), .FEN(FEN[3117]), .op(N8200_t0) );
fim FAN_N8200_1 ( .fault(fault), .net(N8200), .FEN(FEN[3118]), .op(N8200_t1) );
fim FAN_N8204_0 ( .fault(fault), .net(N8204), .FEN(FEN[3119]), .op(N8204_t0) );
fim FAN_N8204_1 ( .fault(fault), .net(N8204), .FEN(FEN[3120]), .op(N8204_t1) );
fim FAN_N8208_0 ( .fault(fault), .net(N8208), .FEN(FEN[3121]), .op(N8208_t0) );
fim FAN_N8208_1 ( .fault(fault), .net(N8208), .FEN(FEN[3122]), .op(N8208_t1) );
fim FAN_N7852_0 ( .fault(fault), .net(N7852), .FEN(FEN[3123]), .op(N7852_t0) );
fim FAN_N7852_1 ( .fault(fault), .net(N7852), .FEN(FEN[3124]), .op(N7852_t1) );
fim FAN_N8114_0 ( .fault(fault), .net(N8114), .FEN(FEN[3125]), .op(N8114_t0) );
fim FAN_N8114_1 ( .fault(fault), .net(N8114), .FEN(FEN[3126]), .op(N8114_t1) );
fim FAN_N7613_0 ( .fault(fault), .net(N7613), .FEN(FEN[3127]), .op(N7613_t0) );
fim FAN_N7613_1 ( .fault(fault), .net(N7613), .FEN(FEN[3128]), .op(N7613_t1) );
fim FAN_N8117_0 ( .fault(fault), .net(N8117), .FEN(FEN[3129]), .op(N8117_t0) );
fim FAN_N8117_1 ( .fault(fault), .net(N8117), .FEN(FEN[3130]), .op(N8117_t1) );
fim FAN_N8131_0 ( .fault(fault), .net(N8131), .FEN(FEN[3131]), .op(N8131_t0) );
fim FAN_N8131_1 ( .fault(fault), .net(N8131), .FEN(FEN[3132]), .op(N8131_t1) );
fim FAN_N8134_0 ( .fault(fault), .net(N8134), .FEN(FEN[3133]), .op(N8134_t0) );
fim FAN_N8134_1 ( .fault(fault), .net(N8134), .FEN(FEN[3134]), .op(N8134_t1) );
fim FAN_N7650_0 ( .fault(fault), .net(N7650), .FEN(FEN[3135]), .op(N7650_t0) );
fim FAN_N7650_1 ( .fault(fault), .net(N7650), .FEN(FEN[3136]), .op(N7650_t1) );
fim FAN_N8146_0 ( .fault(fault), .net(N8146), .FEN(FEN[3137]), .op(N8146_t0) );
fim FAN_N8146_1 ( .fault(fault), .net(N8146), .FEN(FEN[3138]), .op(N8146_t1) );
fim FAN_N8156_0 ( .fault(fault), .net(N8156), .FEN(FEN[3139]), .op(N8156_t0) );
fim FAN_N8156_1 ( .fault(fault), .net(N8156), .FEN(FEN[3140]), .op(N8156_t1) );
fim FAN_N8166_0 ( .fault(fault), .net(N8166), .FEN(FEN[3141]), .op(N8166_t0) );
fim FAN_N8166_1 ( .fault(fault), .net(N8166), .FEN(FEN[3142]), .op(N8166_t1) );
fim FAN_N7659_0 ( .fault(fault), .net(N7659), .FEN(FEN[3143]), .op(N7659_t0) );
fim FAN_N7659_1 ( .fault(fault), .net(N7659), .FEN(FEN[3144]), .op(N7659_t1) );
fim FAN_N8169_0 ( .fault(fault), .net(N8169), .FEN(FEN[3145]), .op(N8169_t0) );
fim FAN_N8169_1 ( .fault(fault), .net(N8169), .FEN(FEN[3146]), .op(N8169_t1) );
fim FAN_N8183_0 ( .fault(fault), .net(N8183), .FEN(FEN[3147]), .op(N8183_t0) );
fim FAN_N8183_1 ( .fault(fault), .net(N8183), .FEN(FEN[3148]), .op(N8183_t1) );
fim FAN_N8186_0 ( .fault(fault), .net(N8186), .FEN(FEN[3149]), .op(N8186_t0) );
fim FAN_N8186_1 ( .fault(fault), .net(N8186), .FEN(FEN[3150]), .op(N8186_t1) );
fim FAN_N8580_0 ( .fault(fault), .net(N8580), .FEN(FEN[3151]), .op(N8580_t0) );
fim FAN_N8580_1 ( .fault(fault), .net(N8580), .FEN(FEN[3152]), .op(N8580_t1) );
fim FAN_N8583_0 ( .fault(fault), .net(N8583), .FEN(FEN[3153]), .op(N8583_t0) );
fim FAN_N8583_1 ( .fault(fault), .net(N8583), .FEN(FEN[3154]), .op(N8583_t1) );
fim FAN_N8586_0 ( .fault(fault), .net(N8586), .FEN(FEN[3155]), .op(N8586_t0) );
fim FAN_N8586_1 ( .fault(fault), .net(N8586), .FEN(FEN[3156]), .op(N8586_t1) );
fim FAN_N8589_0 ( .fault(fault), .net(N8589), .FEN(FEN[3157]), .op(N8589_t0) );
fim FAN_N8589_1 ( .fault(fault), .net(N8589), .FEN(FEN[3158]), .op(N8589_t1) );
fim FAN_N8592_0 ( .fault(fault), .net(N8592), .FEN(FEN[3159]), .op(N8592_t0) );
fim FAN_N8592_1 ( .fault(fault), .net(N8592), .FEN(FEN[3160]), .op(N8592_t1) );
fim FAN_N8595_0 ( .fault(fault), .net(N8595), .FEN(FEN[3161]), .op(N8595_t0) );
fim FAN_N8595_1 ( .fault(fault), .net(N8595), .FEN(FEN[3162]), .op(N8595_t1) );
fim FAN_N8598_0 ( .fault(fault), .net(N8598), .FEN(FEN[3163]), .op(N8598_t0) );
fim FAN_N8598_1 ( .fault(fault), .net(N8598), .FEN(FEN[3164]), .op(N8598_t1) );
fim FAN_N8601_0 ( .fault(fault), .net(N8601), .FEN(FEN[3165]), .op(N8601_t0) );
fim FAN_N8601_1 ( .fault(fault), .net(N8601), .FEN(FEN[3166]), .op(N8601_t1) );
fim FAN_N8604_0 ( .fault(fault), .net(N8604), .FEN(FEN[3167]), .op(N8604_t0) );
fim FAN_N8604_1 ( .fault(fault), .net(N8604), .FEN(FEN[3168]), .op(N8604_t1) );
fim FAN_N8627_0 ( .fault(fault), .net(N8627), .FEN(FEN[3169]), .op(N8627_t0) );
fim FAN_N8627_1 ( .fault(fault), .net(N8627), .FEN(FEN[3170]), .op(N8627_t1) );
fim FAN_N8333_0 ( .fault(fault), .net(N8333), .FEN(FEN[3171]), .op(N8333_t0) );
fim FAN_N8333_1 ( .fault(fault), .net(N8333), .FEN(FEN[3172]), .op(N8333_t1) );
fim FAN_N8333_2 ( .fault(fault), .net(N8333), .FEN(FEN[3173]), .op(N8333_t2) );
fim FAN_N8326_0 ( .fault(fault), .net(N8326), .FEN(FEN[3174]), .op(N8326_t0) );
fim FAN_N8326_1 ( .fault(fault), .net(N8326), .FEN(FEN[3175]), .op(N8326_t1) );
fim FAN_N8326_2 ( .fault(fault), .net(N8326), .FEN(FEN[3176]), .op(N8326_t2) );
fim FAN_N8326_3 ( .fault(fault), .net(N8326), .FEN(FEN[3177]), .op(N8326_t3) );
fim FAN_N8326_4 ( .fault(fault), .net(N8326), .FEN(FEN[3178]), .op(N8326_t4) );
fim FAN_N8326_5 ( .fault(fault), .net(N8326), .FEN(FEN[3179]), .op(N8326_t5) );
fim FAN_N8660_0 ( .fault(fault), .net(N8660), .FEN(FEN[3180]), .op(N8660_t0) );
fim FAN_N8660_1 ( .fault(fault), .net(N8660), .FEN(FEN[3181]), .op(N8660_t1) );
fim FAN_N8663_0 ( .fault(fault), .net(N8663), .FEN(FEN[3182]), .op(N8663_t0) );
fim FAN_N8663_1 ( .fault(fault), .net(N8663), .FEN(FEN[3183]), .op(N8663_t1) );
fim FAN_N8666_0 ( .fault(fault), .net(N8666), .FEN(FEN[3184]), .op(N8666_t0) );
fim FAN_N8666_1 ( .fault(fault), .net(N8666), .FEN(FEN[3185]), .op(N8666_t1) );
fim FAN_N8669_0 ( .fault(fault), .net(N8669), .FEN(FEN[3186]), .op(N8669_t0) );
fim FAN_N8669_1 ( .fault(fault), .net(N8669), .FEN(FEN[3187]), .op(N8669_t1) );
fim FAN_N8672_0 ( .fault(fault), .net(N8672), .FEN(FEN[3188]), .op(N8672_t0) );
fim FAN_N8672_1 ( .fault(fault), .net(N8672), .FEN(FEN[3189]), .op(N8672_t1) );
fim FAN_N8675_0 ( .fault(fault), .net(N8675), .FEN(FEN[3190]), .op(N8675_t0) );
fim FAN_N8675_1 ( .fault(fault), .net(N8675), .FEN(FEN[3191]), .op(N8675_t1) );
fim FAN_N8365_0 ( .fault(fault), .net(N8365), .FEN(FEN[3192]), .op(N8365_t0) );
fim FAN_N8365_1 ( .fault(fault), .net(N8365), .FEN(FEN[3193]), .op(N8365_t1) );
fim FAN_N8365_2 ( .fault(fault), .net(N8365), .FEN(FEN[3194]), .op(N8365_t2) );
fim FAN_N8358_0 ( .fault(fault), .net(N8358), .FEN(FEN[3195]), .op(N8358_t0) );
fim FAN_N8358_1 ( .fault(fault), .net(N8358), .FEN(FEN[3196]), .op(N8358_t1) );
fim FAN_N8358_2 ( .fault(fault), .net(N8358), .FEN(FEN[3197]), .op(N8358_t2) );
fim FAN_N8358_3 ( .fault(fault), .net(N8358), .FEN(FEN[3198]), .op(N8358_t3) );
fim FAN_N8358_4 ( .fault(fault), .net(N8358), .FEN(FEN[3199]), .op(N8358_t4) );
fim FAN_N8358_5 ( .fault(fault), .net(N8358), .FEN(FEN[3200]), .op(N8358_t5) );
fim FAN_N8687_0 ( .fault(fault), .net(N8687), .FEN(FEN[3201]), .op(N8687_t0) );
fim FAN_N8687_1 ( .fault(fault), .net(N8687), .FEN(FEN[3202]), .op(N8687_t1) );
fim FAN_N8699_0 ( .fault(fault), .net(N8699), .FEN(FEN[3203]), .op(N8699_t0) );
fim FAN_N8699_1 ( .fault(fault), .net(N8699), .FEN(FEN[3204]), .op(N8699_t1) );
fim FAN_N8711_0 ( .fault(fault), .net(N8711), .FEN(FEN[3205]), .op(N8711_t0) );
fim FAN_N8711_1 ( .fault(fault), .net(N8711), .FEN(FEN[3206]), .op(N8711_t1) );
fim FAN_N8714_0 ( .fault(fault), .net(N8714), .FEN(FEN[3207]), .op(N8714_t0) );
fim FAN_N8714_1 ( .fault(fault), .net(N8714), .FEN(FEN[3208]), .op(N8714_t1) );
fim FAN_N8727_0 ( .fault(fault), .net(N8727), .FEN(FEN[3209]), .op(N8727_t0) );
fim FAN_N8727_1 ( .fault(fault), .net(N8727), .FEN(FEN[3210]), .op(N8727_t1) );
fim FAN_N8730_0 ( .fault(fault), .net(N8730), .FEN(FEN[3211]), .op(N8730_t0) );
fim FAN_N8730_1 ( .fault(fault), .net(N8730), .FEN(FEN[3212]), .op(N8730_t1) );
fim FAN_N8405_0 ( .fault(fault), .net(N8405), .FEN(FEN[3213]), .op(N8405_t0) );
fim FAN_N8405_1 ( .fault(fault), .net(N8405), .FEN(FEN[3214]), .op(N8405_t1) );
fim FAN_N8405_2 ( .fault(fault), .net(N8405), .FEN(FEN[3215]), .op(N8405_t2) );
fim FAN_N8412_0 ( .fault(fault), .net(N8412), .FEN(FEN[3216]), .op(N8412_t0) );
fim FAN_N8412_1 ( .fault(fault), .net(N8412), .FEN(FEN[3217]), .op(N8412_t1) );
fim FAN_N8430_0 ( .fault(fault), .net(N8430), .FEN(FEN[3218]), .op(N8430_t0) );
fim FAN_N8430_1 ( .fault(fault), .net(N8430), .FEN(FEN[3219]), .op(N8430_t1) );
fim FAN_N8444_0 ( .fault(fault), .net(N8444), .FEN(FEN[3220]), .op(N8444_t0) );
fim FAN_N8444_1 ( .fault(fault), .net(N8444), .FEN(FEN[3221]), .op(N8444_t1) );
fim FAN_N8735_0 ( .fault(fault), .net(N8735), .FEN(FEN[3222]), .op(N8735_t0) );
fim FAN_N8735_1 ( .fault(fault), .net(N8735), .FEN(FEN[3223]), .op(N8735_t1) );
fim FAN_N8738_0 ( .fault(fault), .net(N8738), .FEN(FEN[3224]), .op(N8738_t0) );
fim FAN_N8738_1 ( .fault(fault), .net(N8738), .FEN(FEN[3225]), .op(N8738_t1) );
fim FAN_N8741_0 ( .fault(fault), .net(N8741), .FEN(FEN[3226]), .op(N8741_t0) );
fim FAN_N8741_1 ( .fault(fault), .net(N8741), .FEN(FEN[3227]), .op(N8741_t1) );
fim FAN_N8744_0 ( .fault(fault), .net(N8744), .FEN(FEN[3228]), .op(N8744_t0) );
fim FAN_N8744_1 ( .fault(fault), .net(N8744), .FEN(FEN[3229]), .op(N8744_t1) );
fim FAN_N8747_0 ( .fault(fault), .net(N8747), .FEN(FEN[3230]), .op(N8747_t0) );
fim FAN_N8747_1 ( .fault(fault), .net(N8747), .FEN(FEN[3231]), .op(N8747_t1) );
fim FAN_N8750_0 ( .fault(fault), .net(N8750), .FEN(FEN[3232]), .op(N8750_t0) );
fim FAN_N8750_1 ( .fault(fault), .net(N8750), .FEN(FEN[3233]), .op(N8750_t1) );
fim FAN_N8471_0 ( .fault(fault), .net(N8471), .FEN(FEN[3234]), .op(N8471_t0) );
fim FAN_N8471_1 ( .fault(fault), .net(N8471), .FEN(FEN[3235]), .op(N8471_t1) );
fim FAN_N8474_0 ( .fault(fault), .net(N8474), .FEN(FEN[3236]), .op(N8474_t0) );
fim FAN_N8474_1 ( .fault(fault), .net(N8474), .FEN(FEN[3237]), .op(N8474_t1) );
fim FAN_N8477_0 ( .fault(fault), .net(N8477), .FEN(FEN[3238]), .op(N8477_t0) );
fim FAN_N8477_1 ( .fault(fault), .net(N8477), .FEN(FEN[3239]), .op(N8477_t1) );
fim FAN_N8480_0 ( .fault(fault), .net(N8480), .FEN(FEN[3240]), .op(N8480_t0) );
fim FAN_N8480_1 ( .fault(fault), .net(N8480), .FEN(FEN[3241]), .op(N8480_t1) );
fim FAN_N8460_0 ( .fault(fault), .net(N8460), .FEN(FEN[3242]), .op(N8460_t0) );
fim FAN_N8460_1 ( .fault(fault), .net(N8460), .FEN(FEN[3243]), .op(N8460_t1) );
fim FAN_N8457_0 ( .fault(fault), .net(N8457), .FEN(FEN[3244]), .op(N8457_t0) );
fim FAN_N8457_1 ( .fault(fault), .net(N8457), .FEN(FEN[3245]), .op(N8457_t1) );
fim FAN_N8466_0 ( .fault(fault), .net(N8466), .FEN(FEN[3246]), .op(N8466_t0) );
fim FAN_N8466_1 ( .fault(fault), .net(N8466), .FEN(FEN[3247]), .op(N8466_t1) );
fim FAN_N8463_0 ( .fault(fault), .net(N8463), .FEN(FEN[3248]), .op(N8463_t0) );
fim FAN_N8463_1 ( .fault(fault), .net(N8463), .FEN(FEN[3249]), .op(N8463_t1) );
fim FAN_N8497_0 ( .fault(fault), .net(N8497), .FEN(FEN[3250]), .op(N8497_t0) );
fim FAN_N8497_1 ( .fault(fault), .net(N8497), .FEN(FEN[3251]), .op(N8497_t1) );
fim FAN_N8766_0 ( .fault(fault), .net(N8766), .FEN(FEN[3252]), .op(N8766_t0) );
fim FAN_N8766_1 ( .fault(fault), .net(N8766), .FEN(FEN[3253]), .op(N8766_t1) );
fim FAN_N8778_0 ( .fault(fault), .net(N8778), .FEN(FEN[3254]), .op(N8778_t0) );
fim FAN_N8778_1 ( .fault(fault), .net(N8778), .FEN(FEN[3255]), .op(N8778_t1) );
fim FAN_N8793_0 ( .fault(fault), .net(N8793), .FEN(FEN[3256]), .op(N8793_t0) );
fim FAN_N8793_1 ( .fault(fault), .net(N8793), .FEN(FEN[3257]), .op(N8793_t1) );
fim FAN_N8796_0 ( .fault(fault), .net(N8796), .FEN(FEN[3258]), .op(N8796_t0) );
fim FAN_N8796_1 ( .fault(fault), .net(N8796), .FEN(FEN[3259]), .op(N8796_t1) );
fim FAN_N8485_0 ( .fault(fault), .net(N8485), .FEN(FEN[3260]), .op(N8485_t0) );
fim FAN_N8485_1 ( .fault(fault), .net(N8485), .FEN(FEN[3261]), .op(N8485_t1) );
fim FAN_N8525_0 ( .fault(fault), .net(N8525), .FEN(FEN[3262]), .op(N8525_t0) );
fim FAN_N8525_1 ( .fault(fault), .net(N8525), .FEN(FEN[3263]), .op(N8525_t1) );
fim FAN_N8528_0 ( .fault(fault), .net(N8528), .FEN(FEN[3264]), .op(N8528_t0) );
fim FAN_N8528_1 ( .fault(fault), .net(N8528), .FEN(FEN[3265]), .op(N8528_t1) );
fim FAN_N8531_0 ( .fault(fault), .net(N8531), .FEN(FEN[3266]), .op(N8531_t0) );
fim FAN_N8531_1 ( .fault(fault), .net(N8531), .FEN(FEN[3267]), .op(N8531_t1) );
fim FAN_N8534_0 ( .fault(fault), .net(N8534), .FEN(FEN[3268]), .op(N8534_t0) );
fim FAN_N8534_1 ( .fault(fault), .net(N8534), .FEN(FEN[3269]), .op(N8534_t1) );
fim FAN_N8522_0 ( .fault(fault), .net(N8522), .FEN(FEN[3270]), .op(N8522_t0) );
fim FAN_N8522_1 ( .fault(fault), .net(N8522), .FEN(FEN[3271]), .op(N8522_t1) );
fim FAN_N8519_0 ( .fault(fault), .net(N8519), .FEN(FEN[3272]), .op(N8519_t0) );
fim FAN_N8519_1 ( .fault(fault), .net(N8519), .FEN(FEN[3273]), .op(N8519_t1) );
fim FAN_N7328_0 ( .fault(fault), .net(N7328), .FEN(FEN[3274]), .op(N7328_t0) );
fim FAN_N7328_1 ( .fault(fault), .net(N7328), .FEN(FEN[3275]), .op(N7328_t1) );
fim FAN_N7325_0 ( .fault(fault), .net(N7325), .FEN(FEN[3276]), .op(N7325_t0) );
fim FAN_N7325_1 ( .fault(fault), .net(N7325), .FEN(FEN[3277]), .op(N7325_t1) );
fim FAN_N8541_0 ( .fault(fault), .net(N8541), .FEN(FEN[3278]), .op(N8541_t0) );
fim FAN_N8541_1 ( .fault(fault), .net(N8541), .FEN(FEN[3279]), .op(N8541_t1) );
fim FAN_N8541_2 ( .fault(fault), .net(N8541), .FEN(FEN[3280]), .op(N8541_t2) );
fim FAN_N8548_0 ( .fault(fault), .net(N8548), .FEN(FEN[3281]), .op(N8548_t0) );
fim FAN_N8548_1 ( .fault(fault), .net(N8548), .FEN(FEN[3282]), .op(N8548_t1) );
fim FAN_N89_0 ( .fault(fault), .net(N89), .FEN(FEN[3283]), .op(N89_t0) );
fim FAN_N89_1 ( .fault(fault), .net(N89), .FEN(FEN[3284]), .op(N89_t1) );
fim FAN_N89_2 ( .fault(fault), .net(N89), .FEN(FEN[3285]), .op(N89_t2) );
fim FAN_N89_3 ( .fault(fault), .net(N89), .FEN(FEN[3286]), .op(N89_t3) );
fim FAN_N8811_0 ( .fault(fault), .net(N8811), .FEN(FEN[3287]), .op(N8811_t0) );
fim FAN_N8811_1 ( .fault(fault), .net(N8811), .FEN(FEN[3288]), .op(N8811_t1) );
fim FAN_N8566_0 ( .fault(fault), .net(N8566), .FEN(FEN[3289]), .op(N8566_t0) );
fim FAN_N8566_1 ( .fault(fault), .net(N8566), .FEN(FEN[3290]), .op(N8566_t1) );
fim FAN_N8569_0 ( .fault(fault), .net(N8569), .FEN(FEN[3291]), .op(N8569_t0) );
fim FAN_N8569_1 ( .fault(fault), .net(N8569), .FEN(FEN[3292]), .op(N8569_t1) );
fim FAN_N8572_0 ( .fault(fault), .net(N8572), .FEN(FEN[3293]), .op(N8572_t0) );
fim FAN_N8572_1 ( .fault(fault), .net(N8572), .FEN(FEN[3294]), .op(N8572_t1) );
fim FAN_N8575_0 ( .fault(fault), .net(N8575), .FEN(FEN[3295]), .op(N8575_t0) );
fim FAN_N8575_1 ( .fault(fault), .net(N8575), .FEN(FEN[3296]), .op(N8575_t1) );
fim FAN_N8555_0 ( .fault(fault), .net(N8555), .FEN(FEN[3297]), .op(N8555_t0) );
fim FAN_N8555_1 ( .fault(fault), .net(N8555), .FEN(FEN[3298]), .op(N8555_t1) );
fim FAN_N7384_0 ( .fault(fault), .net(N7384), .FEN(FEN[3299]), .op(N7384_t0) );
fim FAN_N7384_1 ( .fault(fault), .net(N7384), .FEN(FEN[3300]), .op(N7384_t1) );
fim FAN_N8561_0 ( .fault(fault), .net(N8561), .FEN(FEN[3301]), .op(N8561_t0) );
fim FAN_N8561_1 ( .fault(fault), .net(N8561), .FEN(FEN[3302]), .op(N8561_t1) );
fim FAN_N8558_0 ( .fault(fault), .net(N8558), .FEN(FEN[3303]), .op(N8558_t0) );
fim FAN_N8558_1 ( .fault(fault), .net(N8558), .FEN(FEN[3304]), .op(N8558_t1) );
fim FAN_N8678_0 ( .fault(fault), .net(N8678), .FEN(FEN[3305]), .op(N8678_t0) );
fim FAN_N8678_1 ( .fault(fault), .net(N8678), .FEN(FEN[3306]), .op(N8678_t1) );
fim FAN_N8681_0 ( .fault(fault), .net(N8681), .FEN(FEN[3307]), .op(N8681_t0) );
fim FAN_N8681_1 ( .fault(fault), .net(N8681), .FEN(FEN[3308]), .op(N8681_t1) );
fim FAN_N8684_0 ( .fault(fault), .net(N8684), .FEN(FEN[3309]), .op(N8684_t0) );
fim FAN_N8684_1 ( .fault(fault), .net(N8684), .FEN(FEN[3310]), .op(N8684_t1) );
fim FAN_N8690_0 ( .fault(fault), .net(N8690), .FEN(FEN[3311]), .op(N8690_t0) );
fim FAN_N8690_1 ( .fault(fault), .net(N8690), .FEN(FEN[3312]), .op(N8690_t1) );
fim FAN_N8693_0 ( .fault(fault), .net(N8693), .FEN(FEN[3313]), .op(N8693_t0) );
fim FAN_N8693_1 ( .fault(fault), .net(N8693), .FEN(FEN[3314]), .op(N8693_t1) );
fim FAN_N8696_0 ( .fault(fault), .net(N8696), .FEN(FEN[3315]), .op(N8696_t0) );
fim FAN_N8696_1 ( .fault(fault), .net(N8696), .FEN(FEN[3316]), .op(N8696_t1) );
fim FAN_N8702_0 ( .fault(fault), .net(N8702), .FEN(FEN[3317]), .op(N8702_t0) );
fim FAN_N8702_1 ( .fault(fault), .net(N8702), .FEN(FEN[3318]), .op(N8702_t1) );
fim FAN_N8705_0 ( .fault(fault), .net(N8705), .FEN(FEN[3319]), .op(N8705_t0) );
fim FAN_N8705_1 ( .fault(fault), .net(N8705), .FEN(FEN[3320]), .op(N8705_t1) );
fim FAN_N8708_0 ( .fault(fault), .net(N8708), .FEN(FEN[3321]), .op(N8708_t0) );
fim FAN_N8708_1 ( .fault(fault), .net(N8708), .FEN(FEN[3322]), .op(N8708_t1) );
fim FAN_N8724_0 ( .fault(fault), .net(N8724), .FEN(FEN[3323]), .op(N8724_t0) );
fim FAN_N8724_1 ( .fault(fault), .net(N8724), .FEN(FEN[3324]), .op(N8724_t1) );
fim FAN_N8718_0 ( .fault(fault), .net(N8718), .FEN(FEN[3325]), .op(N8718_t0) );
fim FAN_N8718_1 ( .fault(fault), .net(N8718), .FEN(FEN[3326]), .op(N8718_t1) );
fim FAN_N8721_0 ( .fault(fault), .net(N8721), .FEN(FEN[3327]), .op(N8721_t0) );
fim FAN_N8721_1 ( .fault(fault), .net(N8721), .FEN(FEN[3328]), .op(N8721_t1) );
fim FAN_N8757_0 ( .fault(fault), .net(N8757), .FEN(FEN[3329]), .op(N8757_t0) );
fim FAN_N8757_1 ( .fault(fault), .net(N8757), .FEN(FEN[3330]), .op(N8757_t1) );
fim FAN_N8760_0 ( .fault(fault), .net(N8760), .FEN(FEN[3331]), .op(N8760_t0) );
fim FAN_N8760_1 ( .fault(fault), .net(N8760), .FEN(FEN[3332]), .op(N8760_t1) );
fim FAN_N8763_0 ( .fault(fault), .net(N8763), .FEN(FEN[3333]), .op(N8763_t0) );
fim FAN_N8763_1 ( .fault(fault), .net(N8763), .FEN(FEN[3334]), .op(N8763_t1) );
fim FAN_N8769_0 ( .fault(fault), .net(N8769), .FEN(FEN[3335]), .op(N8769_t0) );
fim FAN_N8769_1 ( .fault(fault), .net(N8769), .FEN(FEN[3336]), .op(N8769_t1) );
fim FAN_N8772_0 ( .fault(fault), .net(N8772), .FEN(FEN[3337]), .op(N8772_t0) );
fim FAN_N8772_1 ( .fault(fault), .net(N8772), .FEN(FEN[3338]), .op(N8772_t1) );
fim FAN_N8775_0 ( .fault(fault), .net(N8775), .FEN(FEN[3339]), .op(N8775_t0) );
fim FAN_N8775_1 ( .fault(fault), .net(N8775), .FEN(FEN[3340]), .op(N8775_t1) );
fim FAN_N8781_0 ( .fault(fault), .net(N8781), .FEN(FEN[3341]), .op(N8781_t0) );
fim FAN_N8781_1 ( .fault(fault), .net(N8781), .FEN(FEN[3342]), .op(N8781_t1) );
fim FAN_N8784_0 ( .fault(fault), .net(N8784), .FEN(FEN[3343]), .op(N8784_t0) );
fim FAN_N8784_1 ( .fault(fault), .net(N8784), .FEN(FEN[3344]), .op(N8784_t1) );
fim FAN_N8787_0 ( .fault(fault), .net(N8787), .FEN(FEN[3345]), .op(N8787_t0) );
fim FAN_N8787_1 ( .fault(fault), .net(N8787), .FEN(FEN[3346]), .op(N8787_t1) );
fim FAN_N8790_0 ( .fault(fault), .net(N8790), .FEN(FEN[3347]), .op(N8790_t0) );
fim FAN_N8790_1 ( .fault(fault), .net(N8790), .FEN(FEN[3348]), .op(N8790_t1) );
fim FAN_N8808_0 ( .fault(fault), .net(N8808), .FEN(FEN[3349]), .op(N8808_t0) );
fim FAN_N8808_1 ( .fault(fault), .net(N8808), .FEN(FEN[3350]), .op(N8808_t1) );
fim FAN_N8799_0 ( .fault(fault), .net(N8799), .FEN(FEN[3351]), .op(N8799_t0) );
fim FAN_N8799_1 ( .fault(fault), .net(N8799), .FEN(FEN[3352]), .op(N8799_t1) );
fim FAN_N8802_0 ( .fault(fault), .net(N8802), .FEN(FEN[3353]), .op(N8802_t0) );
fim FAN_N8802_1 ( .fault(fault), .net(N8802), .FEN(FEN[3354]), .op(N8802_t1) );
fim FAN_N8805_0 ( .fault(fault), .net(N8805), .FEN(FEN[3355]), .op(N8805_t0) );
fim FAN_N8805_1 ( .fault(fault), .net(N8805), .FEN(FEN[3356]), .op(N8805_t1) );
fim FAN_N8943_0 ( .fault(fault), .net(N8943), .FEN(FEN[3357]), .op(N8943_t0) );
fim FAN_N8943_1 ( .fault(fault), .net(N8943), .FEN(FEN[3358]), .op(N8943_t1) );
fim FAN_N8943_2 ( .fault(fault), .net(N8943), .FEN(FEN[3359]), .op(N8943_t2) );
fim FAN_N8421_0 ( .fault(fault), .net(N8421), .FEN(FEN[3360]), .op(N8421_t0) );
fim FAN_N8421_1 ( .fault(fault), .net(N8421), .FEN(FEN[3361]), .op(N8421_t1) );
fim FAN_N8421_2 ( .fault(fault), .net(N8421), .FEN(FEN[3362]), .op(N8421_t2) );
fim FAN_N8421_3 ( .fault(fault), .net(N8421), .FEN(FEN[3363]), .op(N8421_t3) );
fim FAN_N8421_4 ( .fault(fault), .net(N8421), .FEN(FEN[3364]), .op(N8421_t4) );
fim FAN_N8421_5 ( .fault(fault), .net(N8421), .FEN(FEN[3365]), .op(N8421_t5) );
fim FAN_N8421_6 ( .fault(fault), .net(N8421), .FEN(FEN[3366]), .op(N8421_t6) );
fim FAN_N8421_7 ( .fault(fault), .net(N8421), .FEN(FEN[3367]), .op(N8421_t7) );
fim FAN_N8857_0 ( .fault(fault), .net(N8857), .FEN(FEN[3368]), .op(N8857_t0) );
fim FAN_N8857_1 ( .fault(fault), .net(N8857), .FEN(FEN[3369]), .op(N8857_t1) );
fim FAN_N8857_2 ( .fault(fault), .net(N8857), .FEN(FEN[3370]), .op(N8857_t2) );
fim FAN_N8871_0 ( .fault(fault), .net(N8871), .FEN(FEN[3371]), .op(N8871_t0) );
fim FAN_N8871_1 ( .fault(fault), .net(N8871), .FEN(FEN[3372]), .op(N8871_t1) );
fim FAN_N8898_0 ( .fault(fault), .net(N8898), .FEN(FEN[3373]), .op(N8898_t0) );
fim FAN_N8898_1 ( .fault(fault), .net(N8898), .FEN(FEN[3374]), .op(N8898_t1) );
fim FAN_N8898_2 ( .fault(fault), .net(N8898), .FEN(FEN[3375]), .op(N8898_t2) );
fim FAN_N8902_0 ( .fault(fault), .net(N8902), .FEN(FEN[3376]), .op(N8902_t0) );
fim FAN_N8902_1 ( .fault(fault), .net(N8902), .FEN(FEN[3377]), .op(N8902_t1) );
fim FAN_N9099_0 ( .fault(fault), .net(N9099), .FEN(FEN[3378]), .op(N9099_t0) );
fim FAN_N9099_1 ( .fault(fault), .net(N9099), .FEN(FEN[3379]), .op(N9099_t1) );
fim FAN_N9103_0 ( .fault(fault), .net(N9103), .FEN(FEN[3380]), .op(N9103_t0) );
fim FAN_N9103_1 ( .fault(fault), .net(N9103), .FEN(FEN[3381]), .op(N9103_t1) );
fim FAN_N9107_0 ( .fault(fault), .net(N9107), .FEN(FEN[3382]), .op(N9107_t0) );
fim FAN_N9107_1 ( .fault(fault), .net(N9107), .FEN(FEN[3383]), .op(N9107_t1) );
fim FAN_N9111_0 ( .fault(fault), .net(N9111), .FEN(FEN[3384]), .op(N9111_t0) );
fim FAN_N9111_1 ( .fault(fault), .net(N9111), .FEN(FEN[3385]), .op(N9111_t1) );
fim FAN_N8920_0 ( .fault(fault), .net(N8920), .FEN(FEN[3386]), .op(N8920_t0) );
fim FAN_N8920_1 ( .fault(fault), .net(N8920), .FEN(FEN[3387]), .op(N8920_t1) );
fim FAN_N8920_2 ( .fault(fault), .net(N8920), .FEN(FEN[3388]), .op(N8920_t2) );
fim FAN_N8927_0 ( .fault(fault), .net(N8927), .FEN(FEN[3389]), .op(N8927_t0) );
fim FAN_N8927_1 ( .fault(fault), .net(N8927), .FEN(FEN[3390]), .op(N8927_t1) );
fim FAN_N8927_2 ( .fault(fault), .net(N8927), .FEN(FEN[3391]), .op(N8927_t2) );
fim FAN_N8950_0 ( .fault(fault), .net(N8950), .FEN(FEN[3392]), .op(N8950_t0) );
fim FAN_N8950_1 ( .fault(fault), .net(N8950), .FEN(FEN[3393]), .op(N8950_t1) );
fim FAN_N8950_2 ( .fault(fault), .net(N8950), .FEN(FEN[3394]), .op(N8950_t2) );
fim FAN_N8956_0 ( .fault(fault), .net(N8956), .FEN(FEN[3395]), .op(N8956_t0) );
fim FAN_N8956_1 ( .fault(fault), .net(N8956), .FEN(FEN[3396]), .op(N8956_t1) );
fim FAN_N8966_0 ( .fault(fault), .net(N8966), .FEN(FEN[3397]), .op(N8966_t0) );
fim FAN_N8966_1 ( .fault(fault), .net(N8966), .FEN(FEN[3398]), .op(N8966_t1) );
fim FAN_N9161_0 ( .fault(fault), .net(N9161), .FEN(FEN[3399]), .op(N9161_t0) );
fim FAN_N9161_1 ( .fault(fault), .net(N9161), .FEN(FEN[3400]), .op(N9161_t1) );
fim FAN_N9165_0 ( .fault(fault), .net(N9165), .FEN(FEN[3401]), .op(N9165_t0) );
fim FAN_N9165_1 ( .fault(fault), .net(N9165), .FEN(FEN[3402]), .op(N9165_t1) );
fim FAN_N9169_0 ( .fault(fault), .net(N9169), .FEN(FEN[3403]), .op(N9169_t0) );
fim FAN_N9169_1 ( .fault(fault), .net(N9169), .FEN(FEN[3404]), .op(N9169_t1) );
fim FAN_N9173_0 ( .fault(fault), .net(N9173), .FEN(FEN[3405]), .op(N9173_t0) );
fim FAN_N9173_1 ( .fault(fault), .net(N9173), .FEN(FEN[3406]), .op(N9173_t1) );
fim FAN_N9001_0 ( .fault(fault), .net(N9001), .FEN(FEN[3407]), .op(N9001_t0) );
fim FAN_N9001_1 ( .fault(fault), .net(N9001), .FEN(FEN[3408]), .op(N9001_t1) );
fim FAN_N9001_2 ( .fault(fault), .net(N9001), .FEN(FEN[3409]), .op(N9001_t2) );
fim FAN_N9029_0 ( .fault(fault), .net(N9029), .FEN(FEN[3410]), .op(N9029_t0) );
fim FAN_N9029_1 ( .fault(fault), .net(N9029), .FEN(FEN[3411]), .op(N9029_t1) );
fim FAN_N9029_2 ( .fault(fault), .net(N9029), .FEN(FEN[3412]), .op(N9029_t2) );
fim FAN_N9035_0 ( .fault(fault), .net(N9035), .FEN(FEN[3413]), .op(N9035_t0) );
fim FAN_N9035_1 ( .fault(fault), .net(N9035), .FEN(FEN[3414]), .op(N9035_t1) );
fim FAN_N9068_0 ( .fault(fault), .net(N9068), .FEN(FEN[3415]), .op(N9068_t0) );
fim FAN_N9068_1 ( .fault(fault), .net(N9068), .FEN(FEN[3416]), .op(N9068_t1) );
fim FAN_N9074_0 ( .fault(fault), .net(N9074), .FEN(FEN[3417]), .op(N9074_t0) );
fim FAN_N9074_1 ( .fault(fault), .net(N9074), .FEN(FEN[3418]), .op(N9074_t1) );
fim FAN_N9079_0 ( .fault(fault), .net(N9079), .FEN(FEN[3419]), .op(N9079_t0) );
fim FAN_N9079_1 ( .fault(fault), .net(N9079), .FEN(FEN[3420]), .op(N9079_t1) );
fim FAN_N9083_0 ( .fault(fault), .net(N9083), .FEN(FEN[3421]), .op(N9083_t0) );
fim FAN_N9083_1 ( .fault(fault), .net(N9083), .FEN(FEN[3422]), .op(N9083_t1) );
fim FAN_N9089_0 ( .fault(fault), .net(N9089), .FEN(FEN[3423]), .op(N9089_t0) );
fim FAN_N9089_1 ( .fault(fault), .net(N9089), .FEN(FEN[3424]), .op(N9089_t1) );
fim FAN_N9095_0 ( .fault(fault), .net(N9095), .FEN(FEN[3425]), .op(N9095_t0) );
fim FAN_N9095_1 ( .fault(fault), .net(N9095), .FEN(FEN[3426]), .op(N9095_t1) );
fim FAN_N8924_0 ( .fault(fault), .net(N8924), .FEN(FEN[3427]), .op(N8924_t0) );
fim FAN_N8924_1 ( .fault(fault), .net(N8924), .FEN(FEN[3428]), .op(N8924_t1) );
fim FAN_N9117_0 ( .fault(fault), .net(N9117), .FEN(FEN[3429]), .op(N9117_t0) );
fim FAN_N9117_1 ( .fault(fault), .net(N9117), .FEN(FEN[3430]), .op(N9117_t1) );
fim FAN_N9127_0 ( .fault(fault), .net(N9127), .FEN(FEN[3431]), .op(N9127_t0) );
fim FAN_N9127_1 ( .fault(fault), .net(N9127), .FEN(FEN[3432]), .op(N9127_t1) );
fim FAN_N8931_0 ( .fault(fault), .net(N8931), .FEN(FEN[3433]), .op(N8931_t0) );
fim FAN_N8931_1 ( .fault(fault), .net(N8931), .FEN(FEN[3434]), .op(N8931_t1) );
fim FAN_N9146_0 ( .fault(fault), .net(N9146), .FEN(FEN[3435]), .op(N9146_t0) );
fim FAN_N9146_1 ( .fault(fault), .net(N9146), .FEN(FEN[3436]), .op(N9146_t1) );
fim FAN_N9149_0 ( .fault(fault), .net(N9149), .FEN(FEN[3437]), .op(N9149_t0) );
fim FAN_N9149_1 ( .fault(fault), .net(N9149), .FEN(FEN[3438]), .op(N9149_t1) );
fim FAN_N8996_0 ( .fault(fault), .net(N8996), .FEN(FEN[3439]), .op(N8996_t0) );
fim FAN_N8996_1 ( .fault(fault), .net(N8996), .FEN(FEN[3440]), .op(N8996_t1) );
fim FAN_N9183_0 ( .fault(fault), .net(N9183), .FEN(FEN[3441]), .op(N9183_t0) );
fim FAN_N9183_1 ( .fault(fault), .net(N9183), .FEN(FEN[3442]), .op(N9183_t1) );
fim FAN_N9193_0 ( .fault(fault), .net(N9193), .FEN(FEN[3443]), .op(N9193_t0) );
fim FAN_N9193_1 ( .fault(fault), .net(N9193), .FEN(FEN[3444]), .op(N9193_t1) );
fim FAN_N9203_0 ( .fault(fault), .net(N9203), .FEN(FEN[3445]), .op(N9203_t0) );
fim FAN_N9203_1 ( .fault(fault), .net(N9203), .FEN(FEN[3446]), .op(N9203_t1) );
fim FAN_N9005_0 ( .fault(fault), .net(N9005), .FEN(FEN[3447]), .op(N9005_t0) );
fim FAN_N9005_1 ( .fault(fault), .net(N9005), .FEN(FEN[3448]), .op(N9005_t1) );
fim FAN_N9206_0 ( .fault(fault), .net(N9206), .FEN(FEN[3449]), .op(N9206_t0) );
fim FAN_N9206_1 ( .fault(fault), .net(N9206), .FEN(FEN[3450]), .op(N9206_t1) );
fim FAN_N9220_0 ( .fault(fault), .net(N9220), .FEN(FEN[3451]), .op(N9220_t0) );
fim FAN_N9220_1 ( .fault(fault), .net(N9220), .FEN(FEN[3452]), .op(N9220_t1) );
fim FAN_N9223_0 ( .fault(fault), .net(N9223), .FEN(FEN[3453]), .op(N9223_t0) );
fim FAN_N9223_1 ( .fault(fault), .net(N9223), .FEN(FEN[3454]), .op(N9223_t1) );
fim FAN_N9268_0 ( .fault(fault), .net(N9268), .FEN(FEN[3455]), .op(N9268_t0) );
fim FAN_N9268_1 ( .fault(fault), .net(N9268), .FEN(FEN[3456]), .op(N9268_t1) );
fim FAN_N8269_0 ( .fault(fault), .net(N8269), .FEN(FEN[3457]), .op(N8269_t0) );
fim FAN_N8269_1 ( .fault(fault), .net(N8269), .FEN(FEN[3458]), .op(N8269_t1) );
fim FAN_N8269_2 ( .fault(fault), .net(N8269), .FEN(FEN[3459]), .op(N8269_t2) );
fim FAN_N8269_3 ( .fault(fault), .net(N8269), .FEN(FEN[3460]), .op(N8269_t3) );
fim FAN_N9408_0 ( .fault(fault), .net(N9408), .FEN(FEN[3461]), .op(N9408_t0) );
fim FAN_N9408_1 ( .fault(fault), .net(N9408), .FEN(FEN[3462]), .op(N9408_t1) );
fim FAN_N9408_2 ( .fault(fault), .net(N9408), .FEN(FEN[3463]), .op(N9408_t2) );
fim FAN_N9332_0 ( .fault(fault), .net(N9332), .FEN(FEN[3464]), .op(N9332_t0) );
fim FAN_N9332_1 ( .fault(fault), .net(N9332), .FEN(FEN[3465]), .op(N9332_t1) );
fim FAN_N9332_2 ( .fault(fault), .net(N9332), .FEN(FEN[3466]), .op(N9332_t2) );
fim FAN_N9332_3 ( .fault(fault), .net(N9332), .FEN(FEN[3467]), .op(N9332_t3) );
fim FAN_N9332_4 ( .fault(fault), .net(N9332), .FEN(FEN[3468]), .op(N9332_t4) );
fim FAN_N9332_5 ( .fault(fault), .net(N9332), .FEN(FEN[3469]), .op(N9332_t5) );
fim FAN_N8394_0 ( .fault(fault), .net(N8394), .FEN(FEN[3470]), .op(N8394_t0) );
fim FAN_N8394_1 ( .fault(fault), .net(N8394), .FEN(FEN[3471]), .op(N8394_t1) );
fim FAN_N8394_2 ( .fault(fault), .net(N8394), .FEN(FEN[3472]), .op(N8394_t2) );
fim FAN_N8394_3 ( .fault(fault), .net(N8394), .FEN(FEN[3473]), .op(N8394_t3) );
fim FAN_N8394_4 ( .fault(fault), .net(N8394), .FEN(FEN[3474]), .op(N8394_t4) );
fim FAN_N8394_5 ( .fault(fault), .net(N8394), .FEN(FEN[3475]), .op(N8394_t5) );
fim FAN_N8394_6 ( .fault(fault), .net(N8394), .FEN(FEN[3476]), .op(N8394_t6) );
fim FAN_N8394_7 ( .fault(fault), .net(N8394), .FEN(FEN[3477]), .op(N8394_t7) );
fim FAN_N8394_8 ( .fault(fault), .net(N8394), .FEN(FEN[3478]), .op(N8394_t8) );
fim FAN_N9265_0 ( .fault(fault), .net(N9265), .FEN(FEN[3479]), .op(N9265_t0) );
fim FAN_N9265_1 ( .fault(fault), .net(N9265), .FEN(FEN[3480]), .op(N9265_t1) );
fim FAN_N8262_0 ( .fault(fault), .net(N8262), .FEN(FEN[3481]), .op(N8262_t0) );
fim FAN_N8262_1 ( .fault(fault), .net(N8262), .FEN(FEN[3482]), .op(N8262_t1) );
fim FAN_N8262_2 ( .fault(fault), .net(N8262), .FEN(FEN[3483]), .op(N8262_t2) );
fim FAN_N8262_3 ( .fault(fault), .net(N8262), .FEN(FEN[3484]), .op(N8262_t3) );
fim FAN_N9423_0 ( .fault(fault), .net(N9423), .FEN(FEN[3485]), .op(N9423_t0) );
fim FAN_N9423_1 ( .fault(fault), .net(N9423), .FEN(FEN[3486]), .op(N9423_t1) );
fim FAN_N9280_0 ( .fault(fault), .net(N9280), .FEN(FEN[3487]), .op(N9280_t0) );
fim FAN_N9280_1 ( .fault(fault), .net(N9280), .FEN(FEN[3488]), .op(N9280_t1) );
fim FAN_N9307_0 ( .fault(fault), .net(N9307), .FEN(FEN[3489]), .op(N9307_t0) );
fim FAN_N9307_1 ( .fault(fault), .net(N9307), .FEN(FEN[3490]), .op(N9307_t1) );
fim FAN_N9307_2 ( .fault(fault), .net(N9307), .FEN(FEN[3491]), .op(N9307_t2) );
fim FAN_N9478_0 ( .fault(fault), .net(N9478), .FEN(FEN[3492]), .op(N9478_t0) );
fim FAN_N9478_1 ( .fault(fault), .net(N9478), .FEN(FEN[3493]), .op(N9478_t1) );
fim FAN_N9485_0 ( .fault(fault), .net(N9485), .FEN(FEN[3494]), .op(N9485_t0) );
fim FAN_N9485_1 ( .fault(fault), .net(N9485), .FEN(FEN[3495]), .op(N9485_t1) );
fim FAN_N9488_0 ( .fault(fault), .net(N9488), .FEN(FEN[3496]), .op(N9488_t0) );
fim FAN_N9488_1 ( .fault(fault), .net(N9488), .FEN(FEN[3497]), .op(N9488_t1) );
fim FAN_N9517_0 ( .fault(fault), .net(N9517), .FEN(FEN[3498]), .op(N9517_t0) );
fim FAN_N9517_1 ( .fault(fault), .net(N9517), .FEN(FEN[3499]), .op(N9517_t1) );
fim FAN_N9520_0 ( .fault(fault), .net(N9520), .FEN(FEN[3500]), .op(N9520_t0) );
fim FAN_N9520_1 ( .fault(fault), .net(N9520), .FEN(FEN[3501]), .op(N9520_t1) );
fim FAN_N9426_0 ( .fault(fault), .net(N9426), .FEN(FEN[3502]), .op(N9426_t0) );
fim FAN_N9426_1 ( .fault(fault), .net(N9426), .FEN(FEN[3503]), .op(N9426_t1) );
fim FAN_N9429_0 ( .fault(fault), .net(N9429), .FEN(FEN[3504]), .op(N9429_t0) );
fim FAN_N9429_1 ( .fault(fault), .net(N9429), .FEN(FEN[3505]), .op(N9429_t1) );
fim FAN_N9462_0 ( .fault(fault), .net(N9462), .FEN(FEN[3506]), .op(N9462_t0) );
fim FAN_N9462_1 ( .fault(fault), .net(N9462), .FEN(FEN[3507]), .op(N9462_t1) );
fim FAN_N9473_0 ( .fault(fault), .net(N9473), .FEN(FEN[3508]), .op(N9473_t0) );
fim FAN_N9473_1 ( .fault(fault), .net(N9473), .FEN(FEN[3509]), .op(N9473_t1) );
fim FAN_N9626_0 ( .fault(fault), .net(N9626), .FEN(FEN[3510]), .op(N9626_t0) );
fim FAN_N9626_1 ( .fault(fault), .net(N9626), .FEN(FEN[3511]), .op(N9626_t1) );
fim FAN_N9629_0 ( .fault(fault), .net(N9629), .FEN(FEN[3512]), .op(N9629_t0) );
fim FAN_N9629_1 ( .fault(fault), .net(N9629), .FEN(FEN[3513]), .op(N9629_t1) );
fim FAN_N9632_0 ( .fault(fault), .net(N9632), .FEN(FEN[3514]), .op(N9632_t0) );
fim FAN_N9632_1 ( .fault(fault), .net(N9632), .FEN(FEN[3515]), .op(N9632_t1) );
fim FAN_N9635_0 ( .fault(fault), .net(N9635), .FEN(FEN[3516]), .op(N9635_t0) );
fim FAN_N9635_1 ( .fault(fault), .net(N9635), .FEN(FEN[3517]), .op(N9635_t1) );
fim FAN_N9543_0 ( .fault(fault), .net(N9543), .FEN(FEN[3518]), .op(N9543_t0) );
fim FAN_N9543_1 ( .fault(fault), .net(N9543), .FEN(FEN[3519]), .op(N9543_t1) );
fim FAN_N9650_0 ( .fault(fault), .net(N9650), .FEN(FEN[3520]), .op(N9650_t0) );
fim FAN_N9650_1 ( .fault(fault), .net(N9650), .FEN(FEN[3521]), .op(N9650_t1) );
fim FAN_N9653_0 ( .fault(fault), .net(N9653), .FEN(FEN[3522]), .op(N9653_t0) );
fim FAN_N9653_1 ( .fault(fault), .net(N9653), .FEN(FEN[3523]), .op(N9653_t1) );
fim FAN_N9656_0 ( .fault(fault), .net(N9656), .FEN(FEN[3524]), .op(N9656_t0) );
fim FAN_N9656_1 ( .fault(fault), .net(N9656), .FEN(FEN[3525]), .op(N9656_t1) );
fim FAN_N9551_0 ( .fault(fault), .net(N9551), .FEN(FEN[3526]), .op(N9551_t0) );
fim FAN_N9551_1 ( .fault(fault), .net(N9551), .FEN(FEN[3527]), .op(N9551_t1) );
fim FAN_N9575_0 ( .fault(fault), .net(N9575), .FEN(FEN[3528]), .op(N9575_t0) );
fim FAN_N9575_1 ( .fault(fault), .net(N9575), .FEN(FEN[3529]), .op(N9575_t1) );
fim FAN_N9575_2 ( .fault(fault), .net(N9575), .FEN(FEN[3530]), .op(N9575_t2) );
fim FAN_N9698_0 ( .fault(fault), .net(N9698), .FEN(FEN[3531]), .op(N9698_t0) );
fim FAN_N9698_1 ( .fault(fault), .net(N9698), .FEN(FEN[3532]), .op(N9698_t1) );
fim FAN_N9702_0 ( .fault(fault), .net(N9702), .FEN(FEN[3533]), .op(N9702_t0) );
fim FAN_N9702_1 ( .fault(fault), .net(N9702), .FEN(FEN[3534]), .op(N9702_t1) );
fim FAN_N9608_0 ( .fault(fault), .net(N9608), .FEN(FEN[3535]), .op(N9608_t0) );
fim FAN_N9608_1 ( .fault(fault), .net(N9608), .FEN(FEN[3536]), .op(N9608_t1) );
fim FAN_N9727_0 ( .fault(fault), .net(N9727), .FEN(FEN[3537]), .op(N9727_t0) );
fim FAN_N9727_1 ( .fault(fault), .net(N9727), .FEN(FEN[3538]), .op(N9727_t1) );
fim FAN_N9642_0 ( .fault(fault), .net(N9642), .FEN(FEN[3539]), .op(N9642_t0) );
fim FAN_N9642_1 ( .fault(fault), .net(N9642), .FEN(FEN[3540]), .op(N9642_t1) );
fim FAN_N9646_0 ( .fault(fault), .net(N9646), .FEN(FEN[3541]), .op(N9646_t0) );
fim FAN_N9646_1 ( .fault(fault), .net(N9646), .FEN(FEN[3542]), .op(N9646_t1) );
fim FAN_N9663_0 ( .fault(fault), .net(N9663), .FEN(FEN[3543]), .op(N9663_t0) );
fim FAN_N9663_1 ( .fault(fault), .net(N9663), .FEN(FEN[3544]), .op(N9663_t1) );
fim FAN_N9667_0 ( .fault(fault), .net(N9667), .FEN(FEN[3545]), .op(N9667_t0) );
fim FAN_N9667_1 ( .fault(fault), .net(N9667), .FEN(FEN[3546]), .op(N9667_t1) );
fim FAN_N9671_0 ( .fault(fault), .net(N9671), .FEN(FEN[3547]), .op(N9671_t0) );
fim FAN_N9671_1 ( .fault(fault), .net(N9671), .FEN(FEN[3548]), .op(N9671_t1) );
fim FAN_N9675_0 ( .fault(fault), .net(N9675), .FEN(FEN[3549]), .op(N9675_t0) );
fim FAN_N9675_1 ( .fault(fault), .net(N9675), .FEN(FEN[3550]), .op(N9675_t1) );
fim FAN_N9679_0 ( .fault(fault), .net(N9679), .FEN(FEN[3551]), .op(N9679_t0) );
fim FAN_N9679_1 ( .fault(fault), .net(N9679), .FEN(FEN[3552]), .op(N9679_t1) );
fim FAN_N9682_0 ( .fault(fault), .net(N9682), .FEN(FEN[3553]), .op(N9682_t0) );
fim FAN_N9682_1 ( .fault(fault), .net(N9682), .FEN(FEN[3554]), .op(N9682_t1) );
fim FAN_N9685_0 ( .fault(fault), .net(N9685), .FEN(FEN[3555]), .op(N9685_t0) );
fim FAN_N9685_1 ( .fault(fault), .net(N9685), .FEN(FEN[3556]), .op(N9685_t1) );
fim FAN_N9692_0 ( .fault(fault), .net(N9692), .FEN(FEN[3557]), .op(N9692_t0) );
fim FAN_N9692_1 ( .fault(fault), .net(N9692), .FEN(FEN[3558]), .op(N9692_t1) );
fim FAN_N9707_0 ( .fault(fault), .net(N9707), .FEN(FEN[3559]), .op(N9707_t0) );
fim FAN_N9707_1 ( .fault(fault), .net(N9707), .FEN(FEN[3560]), .op(N9707_t1) );
fim FAN_N9711_0 ( .fault(fault), .net(N9711), .FEN(FEN[3561]), .op(N9711_t0) );
fim FAN_N9711_1 ( .fault(fault), .net(N9711), .FEN(FEN[3562]), .op(N9711_t1) );
fim FAN_N9717_0 ( .fault(fault), .net(N9717), .FEN(FEN[3563]), .op(N9717_t0) );
fim FAN_N9717_1 ( .fault(fault), .net(N9717), .FEN(FEN[3564]), .op(N9717_t1) );
fim FAN_N9723_0 ( .fault(fault), .net(N9723), .FEN(FEN[3565]), .op(N9723_t0) );
fim FAN_N9723_1 ( .fault(fault), .net(N9723), .FEN(FEN[3566]), .op(N9723_t1) );
fim FAN_N9791_0 ( .fault(fault), .net(N9791), .FEN(FEN[3567]), .op(N9791_t0) );
fim FAN_N9791_1 ( .fault(fault), .net(N9791), .FEN(FEN[3568]), .op(N9791_t1) );
fim FAN_N9791_2 ( .fault(fault), .net(N9791), .FEN(FEN[3569]), .op(N9791_t2) );
fim FAN_N8307_0 ( .fault(fault), .net(N8307), .FEN(FEN[3570]), .op(N8307_t0) );
fim FAN_N8307_1 ( .fault(fault), .net(N8307), .FEN(FEN[3571]), .op(N8307_t1) );
fim FAN_N8307_2 ( .fault(fault), .net(N8307), .FEN(FEN[3572]), .op(N8307_t2) );
fim FAN_N8307_3 ( .fault(fault), .net(N8307), .FEN(FEN[3573]), .op(N8307_t3) );
fim FAN_N8307_4 ( .fault(fault), .net(N8307), .FEN(FEN[3574]), .op(N8307_t4) );
fim FAN_N8307_5 ( .fault(fault), .net(N8307), .FEN(FEN[3575]), .op(N8307_t5) );
fim FAN_N9758_0 ( .fault(fault), .net(N9758), .FEN(FEN[3576]), .op(N9758_t0) );
fim FAN_N9758_1 ( .fault(fault), .net(N9758), .FEN(FEN[3577]), .op(N9758_t1) );
fim FAN_N9758_2 ( .fault(fault), .net(N9758), .FEN(FEN[3578]), .op(N9758_t2) );
fim FAN_N9344_0 ( .fault(fault), .net(N9344), .FEN(FEN[3579]), .op(N9344_t0) );
fim FAN_N9344_1 ( .fault(fault), .net(N9344), .FEN(FEN[3580]), .op(N9344_t1) );
fim FAN_N9344_2 ( .fault(fault), .net(N9344), .FEN(FEN[3581]), .op(N9344_t2) );
fim FAN_N9344_3 ( .fault(fault), .net(N9344), .FEN(FEN[3582]), .op(N9344_t3) );
fim FAN_N9344_4 ( .fault(fault), .net(N9344), .FEN(FEN[3583]), .op(N9344_t4) );
fim FAN_N9344_5 ( .fault(fault), .net(N9344), .FEN(FEN[3584]), .op(N9344_t5) );
fim FAN_N9754_0 ( .fault(fault), .net(N9754), .FEN(FEN[3585]), .op(N9754_t0) );
fim FAN_N9754_1 ( .fault(fault), .net(N9754), .FEN(FEN[3586]), .op(N9754_t1) );
fim FAN_N9754_2 ( .fault(fault), .net(N9754), .FEN(FEN[3587]), .op(N9754_t2) );
fim FAN_N9786_0 ( .fault(fault), .net(N9786), .FEN(FEN[3588]), .op(N9786_t0) );
fim FAN_N9786_1 ( .fault(fault), .net(N9786), .FEN(FEN[3589]), .op(N9786_t1) );
fim FAN_N9786_2 ( .fault(fault), .net(N9786), .FEN(FEN[3590]), .op(N9786_t2) );
fim FAN_N9820_0 ( .fault(fault), .net(N9820), .FEN(FEN[3591]), .op(N9820_t0) );
fim FAN_N9820_1 ( .fault(fault), .net(N9820), .FEN(FEN[3592]), .op(N9820_t1) );
fim FAN_N9820_2 ( .fault(fault), .net(N9820), .FEN(FEN[3593]), .op(N9820_t2) );
fim FAN_N9809_0 ( .fault(fault), .net(N9809), .FEN(FEN[3594]), .op(N9809_t0) );
fim FAN_N9809_1 ( .fault(fault), .net(N9809), .FEN(FEN[3595]), .op(N9809_t1) );
fim FAN_N9809_2 ( .fault(fault), .net(N9809), .FEN(FEN[3596]), .op(N9809_t2) );
fim FAN_N8298_0 ( .fault(fault), .net(N8298), .FEN(FEN[3597]), .op(N8298_t0) );
fim FAN_N8298_1 ( .fault(fault), .net(N8298), .FEN(FEN[3598]), .op(N8298_t1) );
fim FAN_N8298_2 ( .fault(fault), .net(N8298), .FEN(FEN[3599]), .op(N8298_t2) );
fim FAN_N8298_3 ( .fault(fault), .net(N8298), .FEN(FEN[3600]), .op(N8298_t3) );
fim FAN_N8298_4 ( .fault(fault), .net(N8298), .FEN(FEN[3601]), .op(N8298_t4) );
fim FAN_N8298_5 ( .fault(fault), .net(N8298), .FEN(FEN[3602]), .op(N8298_t5) );
fim FAN_N9779_0 ( .fault(fault), .net(N9779), .FEN(FEN[3603]), .op(N9779_t0) );
fim FAN_N9779_1 ( .fault(fault), .net(N9779), .FEN(FEN[3604]), .op(N9779_t1) );
fim FAN_N9779_2 ( .fault(fault), .net(N9779), .FEN(FEN[3605]), .op(N9779_t2) );
fim FAN_N9385_0 ( .fault(fault), .net(N9385), .FEN(FEN[3606]), .op(N9385_t0) );
fim FAN_N9385_1 ( .fault(fault), .net(N9385), .FEN(FEN[3607]), .op(N9385_t1) );
fim FAN_N9385_2 ( .fault(fault), .net(N9385), .FEN(FEN[3608]), .op(N9385_t2) );
fim FAN_N9385_3 ( .fault(fault), .net(N9385), .FEN(FEN[3609]), .op(N9385_t3) );
fim FAN_N9385_4 ( .fault(fault), .net(N9385), .FEN(FEN[3610]), .op(N9385_t4) );
fim FAN_N9385_5 ( .fault(fault), .net(N9385), .FEN(FEN[3611]), .op(N9385_t5) );
fim FAN_N9775_0 ( .fault(fault), .net(N9775), .FEN(FEN[3612]), .op(N9775_t0) );
fim FAN_N9775_1 ( .fault(fault), .net(N9775), .FEN(FEN[3613]), .op(N9775_t1) );
fim FAN_N9775_2 ( .fault(fault), .net(N9775), .FEN(FEN[3614]), .op(N9775_t2) );
fim FAN_N9817_0 ( .fault(fault), .net(N9817), .FEN(FEN[3615]), .op(N9817_t0) );
fim FAN_N9817_1 ( .fault(fault), .net(N9817), .FEN(FEN[3616]), .op(N9817_t1) );
fim FAN_N9339_0 ( .fault(fault), .net(N9339), .FEN(FEN[3617]), .op(N9339_t0) );
fim FAN_N9339_1 ( .fault(fault), .net(N9339), .FEN(FEN[3618]), .op(N9339_t1) );
fim FAN_N9925_0 ( .fault(fault), .net(N9925), .FEN(FEN[3619]), .op(N9925_t0) );
fim FAN_N9925_1 ( .fault(fault), .net(N9925), .FEN(FEN[3620]), .op(N9925_t1) );
fim FAN_N9925_2 ( .fault(fault), .net(N9925), .FEN(FEN[3621]), .op(N9925_t2) );
fim FAN_N9925_3 ( .fault(fault), .net(N9925), .FEN(FEN[3622]), .op(N9925_t3) );
fim FAN_N9925_4 ( .fault(fault), .net(N9925), .FEN(FEN[3623]), .op(N9925_t4) );
fim FAN_N9925_5 ( .fault(fault), .net(N9925), .FEN(FEN[3624]), .op(N9925_t5) );
fim FAN_N9932_0 ( .fault(fault), .net(N9932), .FEN(FEN[3625]), .op(N9932_t0) );
fim FAN_N9932_1 ( .fault(fault), .net(N9932), .FEN(FEN[3626]), .op(N9932_t1) );
fim FAN_N9935_0 ( .fault(fault), .net(N9935), .FEN(FEN[3627]), .op(N9935_t0) );
fim FAN_N9935_1 ( .fault(fault), .net(N9935), .FEN(FEN[3628]), .op(N9935_t1) );
fim FAN_N9983_0 ( .fault(fault), .net(N9983), .FEN(FEN[3629]), .op(N9983_t0) );
fim FAN_N9983_1 ( .fault(fault), .net(N9983), .FEN(FEN[3630]), .op(N9983_t1) );
fim FAN_N9986_0 ( .fault(fault), .net(N9986), .FEN(FEN[3631]), .op(N9986_t0) );
fim FAN_N9986_1 ( .fault(fault), .net(N9986), .FEN(FEN[3632]), .op(N9986_t1) );
fim FAN_N9989_0 ( .fault(fault), .net(N9989), .FEN(FEN[3633]), .op(N9989_t0) );
fim FAN_N9989_1 ( .fault(fault), .net(N9989), .FEN(FEN[3634]), .op(N9989_t1) );
fim FAN_N9992_0 ( .fault(fault), .net(N9992), .FEN(FEN[3635]), .op(N9992_t0) );
fim FAN_N9992_1 ( .fault(fault), .net(N9992), .FEN(FEN[3636]), .op(N9992_t1) );
fim FAN_N9949_0 ( .fault(fault), .net(N9949), .FEN(FEN[3637]), .op(N9949_t0) );
fim FAN_N9949_1 ( .fault(fault), .net(N9949), .FEN(FEN[3638]), .op(N9949_t1) );
fim FAN_N10007_0 ( .fault(fault), .net(N10007), .FEN(FEN[3639]), .op(N10007_t0) );
fim FAN_N10007_1 ( .fault(fault), .net(N10007), .FEN(FEN[3640]), .op(N10007_t1) );
fim FAN_N10010_0 ( .fault(fault), .net(N10010), .FEN(FEN[3641]), .op(N10010_t0) );
fim FAN_N10010_1 ( .fault(fault), .net(N10010), .FEN(FEN[3642]), .op(N10010_t1) );
fim FAN_N9961_0 ( .fault(fault), .net(N9961), .FEN(FEN[3643]), .op(N9961_t0) );
fim FAN_N9961_1 ( .fault(fault), .net(N9961), .FEN(FEN[3644]), .op(N9961_t1) );
fim FAN_N9964_0 ( .fault(fault), .net(N9964), .FEN(FEN[3645]), .op(N9964_t0) );
fim FAN_N9964_1 ( .fault(fault), .net(N9964), .FEN(FEN[3646]), .op(N9964_t1) );
fim FAN_N9979_0 ( .fault(fault), .net(N9979), .FEN(FEN[3647]), .op(N9979_t0) );
fim FAN_N9979_1 ( .fault(fault), .net(N9979), .FEN(FEN[3648]), .op(N9979_t1) );
fim FAN_N9999_0 ( .fault(fault), .net(N9999), .FEN(FEN[3649]), .op(N9999_t0) );
fim FAN_N9999_1 ( .fault(fault), .net(N9999), .FEN(FEN[3650]), .op(N9999_t1) );
fim FAN_N10003_0 ( .fault(fault), .net(N10003), .FEN(FEN[3651]), .op(N10003_t0) );
fim FAN_N10003_1 ( .fault(fault), .net(N10003), .FEN(FEN[3652]), .op(N10003_t1) );
fim FAN_N10070_0 ( .fault(fault), .net(N10070), .FEN(FEN[3653]), .op(N10070_t0) );
fim FAN_N10070_1 ( .fault(fault), .net(N10070), .FEN(FEN[3654]), .op(N10070_t1) );
fim FAN_N10073_0 ( .fault(fault), .net(N10073), .FEN(FEN[3655]), .op(N10073_t0) );
fim FAN_N10073_1 ( .fault(fault), .net(N10073), .FEN(FEN[3656]), .op(N10073_t1) );
fim FAN_N10124_0 ( .fault(fault), .net(N10124), .FEN(FEN[3657]), .op(N10124_t0) );
fim FAN_N10124_1 ( .fault(fault), .net(N10124), .FEN(FEN[3658]), .op(N10124_t1) );
fim FAN_N10124_2 ( .fault(fault), .net(N10124), .FEN(FEN[3659]), .op(N10124_t2) );
fim FAN_N10124_3 ( .fault(fault), .net(N10124), .FEN(FEN[3660]), .op(N10124_t3) );
fim FAN_N10124_4 ( .fault(fault), .net(N10124), .FEN(FEN[3661]), .op(N10124_t4) );
fim FAN_N10116_0 ( .fault(fault), .net(N10116), .FEN(FEN[3662]), .op(N10116_t0) );
fim FAN_N10116_1 ( .fault(fault), .net(N10116), .FEN(FEN[3663]), .op(N10116_t1) );
fim FAN_N10141_0 ( .fault(fault), .net(N10141), .FEN(FEN[3664]), .op(N10141_t0) );
fim FAN_N10141_1 ( .fault(fault), .net(N10141), .FEN(FEN[3665]), .op(N10141_t1) );
fim FAN_N10141_2 ( .fault(fault), .net(N10141), .FEN(FEN[3666]), .op(N10141_t2) );
fim FAN_N10141_3 ( .fault(fault), .net(N10141), .FEN(FEN[3667]), .op(N10141_t3) );
fim FAN_N10141_4 ( .fault(fault), .net(N10141), .FEN(FEN[3668]), .op(N10141_t4) );
fim FAN_N10141_5 ( .fault(fault), .net(N10141), .FEN(FEN[3669]), .op(N10141_t5) );
fim FAN_N10119_0 ( .fault(fault), .net(N10119), .FEN(FEN[3670]), .op(N10119_t0) );
fim FAN_N10119_1 ( .fault(fault), .net(N10119), .FEN(FEN[3671]), .op(N10119_t1) );
fim FAN_N10119_2 ( .fault(fault), .net(N10119), .FEN(FEN[3672]), .op(N10119_t2) );
fim FAN_N10119_3 ( .fault(fault), .net(N10119), .FEN(FEN[3673]), .op(N10119_t3) );
fim FAN_N10148_0 ( .fault(fault), .net(N10148), .FEN(FEN[3674]), .op(N10148_t0) );
fim FAN_N10148_1 ( .fault(fault), .net(N10148), .FEN(FEN[3675]), .op(N10148_t1) );
fim FAN_N10148_2 ( .fault(fault), .net(N10148), .FEN(FEN[3676]), .op(N10148_t2) );
fim FAN_N10148_3 ( .fault(fault), .net(N10148), .FEN(FEN[3677]), .op(N10148_t3) );
fim FAN_N10148_4 ( .fault(fault), .net(N10148), .FEN(FEN[3678]), .op(N10148_t4) );
fim FAN_N10148_5 ( .fault(fault), .net(N10148), .FEN(FEN[3679]), .op(N10148_t5) );
fim FAN_N10170_0 ( .fault(fault), .net(N10170), .FEN(FEN[3680]), .op(N10170_t0) );
fim FAN_N10170_1 ( .fault(fault), .net(N10170), .FEN(FEN[3681]), .op(N10170_t1) );
fim FAN_N10173_0 ( .fault(fault), .net(N10173), .FEN(FEN[3682]), .op(N10173_t0) );
fim FAN_N10173_1 ( .fault(fault), .net(N10173), .FEN(FEN[3683]), .op(N10173_t1) );
fim FAN_N10180_0 ( .fault(fault), .net(N10180), .FEN(FEN[3684]), .op(N10180_t0) );
fim FAN_N10180_1 ( .fault(fault), .net(N10180), .FEN(FEN[3685]), .op(N10180_t1) );
fim FAN_N10183_0 ( .fault(fault), .net(N10183), .FEN(FEN[3686]), .op(N10183_t0) );
fim FAN_N10183_1 ( .fault(fault), .net(N10183), .FEN(FEN[3687]), .op(N10183_t1) );
fim FAN_N10186_0 ( .fault(fault), .net(N10186), .FEN(FEN[3688]), .op(N10186_t0) );
fim FAN_N10186_1 ( .fault(fault), .net(N10186), .FEN(FEN[3689]), .op(N10186_t1) );
fim FAN_N10189_0 ( .fault(fault), .net(N10189), .FEN(FEN[3690]), .op(N10189_t0) );
fim FAN_N10189_1 ( .fault(fault), .net(N10189), .FEN(FEN[3691]), .op(N10189_t1) );
fim FAN_N10192_0 ( .fault(fault), .net(N10192), .FEN(FEN[3692]), .op(N10192_t0) );
fim FAN_N10192_1 ( .fault(fault), .net(N10192), .FEN(FEN[3693]), .op(N10192_t1) );
fim FAN_N10197_0 ( .fault(fault), .net(N10197), .FEN(FEN[3694]), .op(N10197_t0) );
fim FAN_N10197_1 ( .fault(fault), .net(N10197), .FEN(FEN[3695]), .op(N10197_t1) );
fim FAN_N10200_0 ( .fault(fault), .net(N10200), .FEN(FEN[3696]), .op(N10200_t0) );
fim FAN_N10200_1 ( .fault(fault), .net(N10200), .FEN(FEN[3697]), .op(N10200_t1) );
fim FAN_N10296_0 ( .fault(fault), .net(N10296), .FEN(FEN[3698]), .op(N10296_t0) );
fim FAN_N10296_1 ( .fault(fault), .net(N10296), .FEN(FEN[3699]), .op(N10296_t1) );
fim FAN_N10308_0 ( .fault(fault), .net(N10308), .FEN(FEN[3700]), .op(N10308_t0) );
fim FAN_N10308_1 ( .fault(fault), .net(N10308), .FEN(FEN[3701]), .op(N10308_t1) );
fim FAN_N10311_0 ( .fault(fault), .net(N10311), .FEN(FEN[3702]), .op(N10311_t0) );
fim FAN_N10311_1 ( .fault(fault), .net(N10311), .FEN(FEN[3703]), .op(N10311_t1) );
fim FAN_N10273_0 ( .fault(fault), .net(N10273), .FEN(FEN[3704]), .op(N10273_t0) );
fim FAN_N10273_1 ( .fault(fault), .net(N10273), .FEN(FEN[3705]), .op(N10273_t1) );
fim FAN_N10273_2 ( .fault(fault), .net(N10273), .FEN(FEN[3706]), .op(N10273_t2) );
fim FAN_N10273_3 ( .fault(fault), .net(N10273), .FEN(FEN[3707]), .op(N10273_t3) );
fim FAN_N10301_0 ( .fault(fault), .net(N10301), .FEN(FEN[3708]), .op(N10301_t0) );
fim FAN_N10301_1 ( .fault(fault), .net(N10301), .FEN(FEN[3709]), .op(N10301_t1) );
fim FAN_N10301_2 ( .fault(fault), .net(N10301), .FEN(FEN[3710]), .op(N10301_t2) );
fim FAN_N10301_3 ( .fault(fault), .net(N10301), .FEN(FEN[3711]), .op(N10301_t3) );
fim FAN_N10318_0 ( .fault(fault), .net(N10318), .FEN(FEN[3712]), .op(N10318_t0) );
fim FAN_N10318_1 ( .fault(fault), .net(N10318), .FEN(FEN[3713]), .op(N10318_t1) );
fim FAN_N10321_0 ( .fault(fault), .net(N10321), .FEN(FEN[3714]), .op(N10321_t0) );
fim FAN_N10321_1 ( .fault(fault), .net(N10321), .FEN(FEN[3715]), .op(N10321_t1) );
fim FAN_N10334_0 ( .fault(fault), .net(N10334), .FEN(FEN[3716]), .op(N10334_t0) );
fim FAN_N10334_1 ( .fault(fault), .net(N10334), .FEN(FEN[3717]), .op(N10334_t1) );
fim FAN_N10341_0 ( .fault(fault), .net(N10341), .FEN(FEN[3718]), .op(N10341_t0) );
fim FAN_N10341_1 ( .fault(fault), .net(N10341), .FEN(FEN[3719]), .op(N10341_t1) );
fim FAN_N10344_0 ( .fault(fault), .net(N10344), .FEN(FEN[3720]), .op(N10344_t0) );
fim FAN_N10344_1 ( .fault(fault), .net(N10344), .FEN(FEN[3721]), .op(N10344_t1) );
fim FAN_N10391_0 ( .fault(fault), .net(N10391), .FEN(FEN[3722]), .op(N10391_t0) );
fim FAN_N10391_1 ( .fault(fault), .net(N10391), .FEN(FEN[3723]), .op(N10391_t1) );
fim FAN_N10367_0 ( .fault(fault), .net(N10367), .FEN(FEN[3724]), .op(N10367_t0) );
fim FAN_N10367_1 ( .fault(fault), .net(N10367), .FEN(FEN[3725]), .op(N10367_t1) );
fim FAN_N10367_2 ( .fault(fault), .net(N10367), .FEN(FEN[3726]), .op(N10367_t2) );
fim FAN_N10367_3 ( .fault(fault), .net(N10367), .FEN(FEN[3727]), .op(N10367_t3) );
fim FAN_N10354_0 ( .fault(fault), .net(N10354), .FEN(FEN[3728]), .op(N10354_t0) );
fim FAN_N10354_1 ( .fault(fault), .net(N10354), .FEN(FEN[3729]), .op(N10354_t1) );
fim FAN_N10375_0 ( .fault(fault), .net(N10375), .FEN(FEN[3730]), .op(N10375_t0) );
fim FAN_N10375_1 ( .fault(fault), .net(N10375), .FEN(FEN[3731]), .op(N10375_t1) );
fim FAN_N10375_2 ( .fault(fault), .net(N10375), .FEN(FEN[3732]), .op(N10375_t2) );
fim FAN_N10375_3 ( .fault(fault), .net(N10375), .FEN(FEN[3733]), .op(N10375_t3) );
fim FAN_N10375_4 ( .fault(fault), .net(N10375), .FEN(FEN[3734]), .op(N10375_t4) );
fim FAN_N10406_0 ( .fault(fault), .net(N10406), .FEN(FEN[3735]), .op(N10406_t0) );
fim FAN_N10406_1 ( .fault(fault), .net(N10406), .FEN(FEN[3736]), .op(N10406_t1) );
fim FAN_N10409_0 ( .fault(fault), .net(N10409), .FEN(FEN[3737]), .op(N10409_t0) );
fim FAN_N10409_1 ( .fault(fault), .net(N10409), .FEN(FEN[3738]), .op(N10409_t1) );
fim FAN_N10412_0 ( .fault(fault), .net(N10412), .FEN(FEN[3739]), .op(N10412_t0) );
fim FAN_N10412_1 ( .fault(fault), .net(N10412), .FEN(FEN[3740]), .op(N10412_t1) );
fim FAN_N10415_0 ( .fault(fault), .net(N10415), .FEN(FEN[3741]), .op(N10415_t0) );
fim FAN_N10415_1 ( .fault(fault), .net(N10415), .FEN(FEN[3742]), .op(N10415_t1) );
fim FAN_N10419_0 ( .fault(fault), .net(N10419), .FEN(FEN[3743]), .op(N10419_t0) );
fim FAN_N10419_1 ( .fault(fault), .net(N10419), .FEN(FEN[3744]), .op(N10419_t1) );
fim FAN_N10422_0 ( .fault(fault), .net(N10422), .FEN(FEN[3745]), .op(N10422_t0) );
fim FAN_N10422_1 ( .fault(fault), .net(N10422), .FEN(FEN[3746]), .op(N10422_t1) );
fim FAN_N10425_0 ( .fault(fault), .net(N10425), .FEN(FEN[3747]), .op(N10425_t0) );
fim FAN_N10425_1 ( .fault(fault), .net(N10425), .FEN(FEN[3748]), .op(N10425_t1) );
fim FAN_N10428_0 ( .fault(fault), .net(N10428), .FEN(FEN[3749]), .op(N10428_t0) );
fim FAN_N10428_1 ( .fault(fault), .net(N10428), .FEN(FEN[3750]), .op(N10428_t1) );
fim FAN_N10399_0 ( .fault(fault), .net(N10399), .FEN(FEN[3751]), .op(N10399_t0) );
fim FAN_N10399_1 ( .fault(fault), .net(N10399), .FEN(FEN[3752]), .op(N10399_t1) );
fim FAN_N10402_0 ( .fault(fault), .net(N10402), .FEN(FEN[3753]), .op(N10402_t0) );
fim FAN_N10402_1 ( .fault(fault), .net(N10402), .FEN(FEN[3754]), .op(N10402_t1) );
fim FAN_N10388_0 ( .fault(fault), .net(N10388), .FEN(FEN[3755]), .op(N10388_t0) );
fim FAN_N10388_1 ( .fault(fault), .net(N10388), .FEN(FEN[3756]), .op(N10388_t1) );
fim FAN_N10360_0 ( .fault(fault), .net(N10360), .FEN(FEN[3757]), .op(N10360_t0) );
fim FAN_N10360_1 ( .fault(fault), .net(N10360), .FEN(FEN[3758]), .op(N10360_t1) );
fim FAN_N10357_0 ( .fault(fault), .net(N10357), .FEN(FEN[3759]), .op(N10357_t0) );
fim FAN_N10357_1 ( .fault(fault), .net(N10357), .FEN(FEN[3760]), .op(N10357_t1) );
fim FAN_N10381_0 ( .fault(fault), .net(N10381), .FEN(FEN[3761]), .op(N10381_t0) );
fim FAN_N10381_1 ( .fault(fault), .net(N10381), .FEN(FEN[3762]), .op(N10381_t1) );
fim FAN_N10381_2 ( .fault(fault), .net(N10381), .FEN(FEN[3763]), .op(N10381_t2) );
fim FAN_N10381_3 ( .fault(fault), .net(N10381), .FEN(FEN[3764]), .op(N10381_t3) );
fim FAN_N10381_4 ( .fault(fault), .net(N10381), .FEN(FEN[3765]), .op(N10381_t4) );
fim FAN_N10381_5 ( .fault(fault), .net(N10381), .FEN(FEN[3766]), .op(N10381_t5) );
fim FAN_N10479_0 ( .fault(fault), .net(N10479), .FEN(FEN[3767]), .op(N10479_t0) );
fim FAN_N10479_1 ( .fault(fault), .net(N10479), .FEN(FEN[3768]), .op(N10479_t1) );
fim FAN_N10479_2 ( .fault(fault), .net(N10479), .FEN(FEN[3769]), .op(N10479_t2) );
fim FAN_N10509_0 ( .fault(fault), .net(N10509), .FEN(FEN[3770]), .op(N10509_t0) );
fim FAN_N10509_1 ( .fault(fault), .net(N10509), .FEN(FEN[3771]), .op(N10509_t1) );
fim FAN_N10512_0 ( .fault(fault), .net(N10512), .FEN(FEN[3772]), .op(N10512_t0) );
fim FAN_N10512_1 ( .fault(fault), .net(N10512), .FEN(FEN[3773]), .op(N10512_t1) );
fim FAN_N10519_0 ( .fault(fault), .net(N10519), .FEN(FEN[3774]), .op(N10519_t0) );
fim FAN_N10519_1 ( .fault(fault), .net(N10519), .FEN(FEN[3775]), .op(N10519_t1) );
fim FAN_N10522_0 ( .fault(fault), .net(N10522), .FEN(FEN[3776]), .op(N10522_t0) );
fim FAN_N10522_1 ( .fault(fault), .net(N10522), .FEN(FEN[3777]), .op(N10522_t1) );
fim FAN_N10525_0 ( .fault(fault), .net(N10525), .FEN(FEN[3778]), .op(N10525_t0) );
fim FAN_N10525_1 ( .fault(fault), .net(N10525), .FEN(FEN[3779]), .op(N10525_t1) );
fim FAN_N10528_0 ( .fault(fault), .net(N10528), .FEN(FEN[3780]), .op(N10528_t0) );
fim FAN_N10528_1 ( .fault(fault), .net(N10528), .FEN(FEN[3781]), .op(N10528_t1) );
fim FAN_N10531_0 ( .fault(fault), .net(N10531), .FEN(FEN[3782]), .op(N10531_t0) );
fim FAN_N10531_1 ( .fault(fault), .net(N10531), .FEN(FEN[3783]), .op(N10531_t1) );
fim FAN_N10536_0 ( .fault(fault), .net(N10536), .FEN(FEN[3784]), .op(N10536_t0) );
fim FAN_N10536_1 ( .fault(fault), .net(N10536), .FEN(FEN[3785]), .op(N10536_t1) );
fim FAN_N10539_0 ( .fault(fault), .net(N10539), .FEN(FEN[3786]), .op(N10539_t0) );
fim FAN_N10539_1 ( .fault(fault), .net(N10539), .FEN(FEN[3787]), .op(N10539_t1) );
fim FAN_N10583_0 ( .fault(fault), .net(N10583), .FEN(FEN[3788]), .op(N10583_t0) );
fim FAN_N10583_1 ( .fault(fault), .net(N10583), .FEN(FEN[3789]), .op(N10583_t1) );
fim FAN_N10583_2 ( .fault(fault), .net(N10583), .FEN(FEN[3790]), .op(N10583_t2) );
fim FAN_N10589_0 ( .fault(fault), .net(N10589), .FEN(FEN[3791]), .op(N10589_t0) );
fim FAN_N10589_1 ( .fault(fault), .net(N10589), .FEN(FEN[3792]), .op(N10589_t1) );
fim FAN_N10589_2 ( .fault(fault), .net(N10589), .FEN(FEN[3793]), .op(N10589_t2) );
fim FAN_N10589_3 ( .fault(fault), .net(N10589), .FEN(FEN[3794]), .op(N10589_t3) );
fim FAN_N10602_0 ( .fault(fault), .net(N10602), .FEN(FEN[3795]), .op(N10602_t0) );
fim FAN_N10602_1 ( .fault(fault), .net(N10602), .FEN(FEN[3796]), .op(N10602_t1) );
fim FAN_N10652_0 ( .fault(fault), .net(N10652), .FEN(FEN[3797]), .op(N10652_t0) );
fim FAN_N10652_1 ( .fault(fault), .net(N10652), .FEN(FEN[3798]), .op(N10652_t1) );
fim FAN_N10652_2 ( .fault(fault), .net(N10652), .FEN(FEN[3799]), .op(N10652_t2) );
fim FAN_N10652_3 ( .fault(fault), .net(N10652), .FEN(FEN[3800]), .op(N10652_t3) );
fim FAN_N10652_4 ( .fault(fault), .net(N10652), .FEN(FEN[3801]), .op(N10652_t4) );
fim FAN_N10659_0 ( .fault(fault), .net(N10659), .FEN(FEN[3802]), .op(N10659_t0) );
fim FAN_N10659_1 ( .fault(fault), .net(N10659), .FEN(FEN[3803]), .op(N10659_t1) );
fim FAN_N10662_0 ( .fault(fault), .net(N10662), .FEN(FEN[3804]), .op(N10662_t0) );
fim FAN_N10662_1 ( .fault(fault), .net(N10662), .FEN(FEN[3805]), .op(N10662_t1) );
fim FAN_N10665_0 ( .fault(fault), .net(N10665), .FEN(FEN[3806]), .op(N10665_t0) );
fim FAN_N10665_1 ( .fault(fault), .net(N10665), .FEN(FEN[3807]), .op(N10665_t1) );
fim FAN_N10668_0 ( .fault(fault), .net(N10668), .FEN(FEN[3808]), .op(N10668_t0) );
fim FAN_N10668_1 ( .fault(fault), .net(N10668), .FEN(FEN[3809]), .op(N10668_t1) );
fim FAN_N10675_0 ( .fault(fault), .net(N10675), .FEN(FEN[3810]), .op(N10675_t0) );
fim FAN_N10675_1 ( .fault(fault), .net(N10675), .FEN(FEN[3811]), .op(N10675_t1) );
fim FAN_N10678_0 ( .fault(fault), .net(N10678), .FEN(FEN[3812]), .op(N10678_t0) );
fim FAN_N10678_1 ( .fault(fault), .net(N10678), .FEN(FEN[3813]), .op(N10678_t1) );
fim FAN_N10691_0 ( .fault(fault), .net(N10691), .FEN(FEN[3814]), .op(N10691_t0) );
fim FAN_N10691_1 ( .fault(fault), .net(N10691), .FEN(FEN[3815]), .op(N10691_t1) );
fim FAN_N10698_0 ( .fault(fault), .net(N10698), .FEN(FEN[3816]), .op(N10698_t0) );
fim FAN_N10698_1 ( .fault(fault), .net(N10698), .FEN(FEN[3817]), .op(N10698_t1) );
fim FAN_N10701_0 ( .fault(fault), .net(N10701), .FEN(FEN[3818]), .op(N10701_t0) );
fim FAN_N10701_1 ( .fault(fault), .net(N10701), .FEN(FEN[3819]), .op(N10701_t1) );
fim FAN_N10739_0 ( .fault(fault), .net(N10739), .FEN(FEN[3820]), .op(N10739_t0) );
fim FAN_N10739_1 ( .fault(fault), .net(N10739), .FEN(FEN[3821]), .op(N10739_t1) );
fim FAN_N10778_0 ( .fault(fault), .net(N10778), .FEN(FEN[3822]), .op(N10778_t0) );
fim FAN_N10778_1 ( .fault(fault), .net(N10778), .FEN(FEN[3823]), .op(N10778_t1) );
fim FAN_N10781_0 ( .fault(fault), .net(N10781), .FEN(FEN[3824]), .op(N10781_t0) );
fim FAN_N10781_1 ( .fault(fault), .net(N10781), .FEN(FEN[3825]), .op(N10781_t1) );
fim FAN_N10784_0 ( .fault(fault), .net(N10784), .FEN(FEN[3826]), .op(N10784_t0) );
fim FAN_N10784_1 ( .fault(fault), .net(N10784), .FEN(FEN[3827]), .op(N10784_t1) );
fim FAN_N10784_2 ( .fault(fault), .net(N10784), .FEN(FEN[3828]), .op(N10784_t2) );
fim FAN_N10784_3 ( .fault(fault), .net(N10784), .FEN(FEN[3829]), .op(N10784_t3) );
fim FAN_N10789_0 ( .fault(fault), .net(N10789), .FEN(FEN[3830]), .op(N10789_t0) );
fim FAN_N10789_1 ( .fault(fault), .net(N10789), .FEN(FEN[3831]), .op(N10789_t1) );
fim FAN_N10792_0 ( .fault(fault), .net(N10792), .FEN(FEN[3832]), .op(N10792_t0) );
fim FAN_N10792_1 ( .fault(fault), .net(N10792), .FEN(FEN[3833]), .op(N10792_t1) );
fim FAN_N10800_0 ( .fault(fault), .net(N10800), .FEN(FEN[3834]), .op(N10800_t0) );
fim FAN_N10800_1 ( .fault(fault), .net(N10800), .FEN(FEN[3835]), .op(N10800_t1) );
fim FAN_N10803_0 ( .fault(fault), .net(N10803), .FEN(FEN[3836]), .op(N10803_t0) );
fim FAN_N10803_1 ( .fault(fault), .net(N10803), .FEN(FEN[3837]), .op(N10803_t1) );
fim FAN_N10806_0 ( .fault(fault), .net(N10806), .FEN(FEN[3838]), .op(N10806_t0) );
fim FAN_N10806_1 ( .fault(fault), .net(N10806), .FEN(FEN[3839]), .op(N10806_t1) );
fim FAN_N10809_0 ( .fault(fault), .net(N10809), .FEN(FEN[3840]), .op(N10809_t0) );
fim FAN_N10809_1 ( .fault(fault), .net(N10809), .FEN(FEN[3841]), .op(N10809_t1) );
fim FAN_N10812_0 ( .fault(fault), .net(N10812), .FEN(FEN[3842]), .op(N10812_t0) );
fim FAN_N10812_1 ( .fault(fault), .net(N10812), .FEN(FEN[3843]), .op(N10812_t1) );
fim FAN_N10817_0 ( .fault(fault), .net(N10817), .FEN(FEN[3844]), .op(N10817_t0) );
fim FAN_N10817_1 ( .fault(fault), .net(N10817), .FEN(FEN[3845]), .op(N10817_t1) );
fim FAN_N10820_0 ( .fault(fault), .net(N10820), .FEN(FEN[3846]), .op(N10820_t0) );
fim FAN_N10820_1 ( .fault(fault), .net(N10820), .FEN(FEN[3847]), .op(N10820_t1) );
fim FAN_N10876_0 ( .fault(fault), .net(N10876), .FEN(FEN[3848]), .op(N10876_t0) );
fim FAN_N10876_1 ( .fault(fault), .net(N10876), .FEN(FEN[3849]), .op(N10876_t1) );
fim FAN_N10879_0 ( .fault(fault), .net(N10879), .FEN(FEN[3850]), .op(N10879_t0) );
fim FAN_N10879_1 ( .fault(fault), .net(N10879), .FEN(FEN[3851]), .op(N10879_t1) );
fim FAN_N10892_0 ( .fault(fault), .net(N10892), .FEN(FEN[3852]), .op(N10892_t0) );
fim FAN_N10892_1 ( .fault(fault), .net(N10892), .FEN(FEN[3853]), .op(N10892_t1) );
fim FAN_N10899_0 ( .fault(fault), .net(N10899), .FEN(FEN[3854]), .op(N10899_t0) );
fim FAN_N10899_1 ( .fault(fault), .net(N10899), .FEN(FEN[3855]), .op(N10899_t1) );
fim FAN_N10902_0 ( .fault(fault), .net(N10902), .FEN(FEN[3856]), .op(N10902_t0) );
fim FAN_N10902_1 ( .fault(fault), .net(N10902), .FEN(FEN[3857]), .op(N10902_t1) );
fim FAN_N10928_0 ( .fault(fault), .net(N10928), .FEN(FEN[3858]), .op(N10928_t0) );
fim FAN_N10928_1 ( .fault(fault), .net(N10928), .FEN(FEN[3859]), .op(N10928_t1) );
fim FAN_N10931_0 ( .fault(fault), .net(N10931), .FEN(FEN[3860]), .op(N10931_t0) );
fim FAN_N10931_1 ( .fault(fault), .net(N10931), .FEN(FEN[3861]), .op(N10931_t1) );
fim FAN_N10938_0 ( .fault(fault), .net(N10938), .FEN(FEN[3862]), .op(N10938_t0) );
fim FAN_N10938_1 ( .fault(fault), .net(N10938), .FEN(FEN[3863]), .op(N10938_t1) );
fim FAN_N10941_0 ( .fault(fault), .net(N10941), .FEN(FEN[3864]), .op(N10941_t0) );
fim FAN_N10941_1 ( .fault(fault), .net(N10941), .FEN(FEN[3865]), .op(N10941_t1) );
fim FAN_N10944_0 ( .fault(fault), .net(N10944), .FEN(FEN[3866]), .op(N10944_t0) );
fim FAN_N10944_1 ( .fault(fault), .net(N10944), .FEN(FEN[3867]), .op(N10944_t1) );
fim FAN_N10947_0 ( .fault(fault), .net(N10947), .FEN(FEN[3868]), .op(N10947_t0) );
fim FAN_N10947_1 ( .fault(fault), .net(N10947), .FEN(FEN[3869]), .op(N10947_t1) );
fim FAN_N10950_0 ( .fault(fault), .net(N10950), .FEN(FEN[3870]), .op(N10950_t0) );
fim FAN_N10950_1 ( .fault(fault), .net(N10950), .FEN(FEN[3871]), .op(N10950_t1) );
fim FAN_N10955_0 ( .fault(fault), .net(N10955), .FEN(FEN[3872]), .op(N10955_t0) );
fim FAN_N10955_1 ( .fault(fault), .net(N10955), .FEN(FEN[3873]), .op(N10955_t1) );
fim FAN_N10958_0 ( .fault(fault), .net(N10958), .FEN(FEN[3874]), .op(N10958_t0) );
fim FAN_N10958_1 ( .fault(fault), .net(N10958), .FEN(FEN[3875]), .op(N10958_t1) );
fim FAN_N10992_0 ( .fault(fault), .net(N10992), .FEN(FEN[3876]), .op(N10992_t0) );
fim FAN_N10992_1 ( .fault(fault), .net(N10992), .FEN(FEN[3877]), .op(N10992_t1) );
fim FAN_N10995_0 ( .fault(fault), .net(N10995), .FEN(FEN[3878]), .op(N10995_t0) );
fim FAN_N10995_1 ( .fault(fault), .net(N10995), .FEN(FEN[3879]), .op(N10995_t1) );
fim FAN_N11008_0 ( .fault(fault), .net(N11008), .FEN(FEN[3880]), .op(N11008_t0) );
fim FAN_N11008_1 ( .fault(fault), .net(N11008), .FEN(FEN[3881]), .op(N11008_t1) );
fim FAN_N11015_0 ( .fault(fault), .net(N11015), .FEN(FEN[3882]), .op(N11015_t0) );
fim FAN_N11015_1 ( .fault(fault), .net(N11015), .FEN(FEN[3883]), .op(N11015_t1) );
fim FAN_N11018_0 ( .fault(fault), .net(N11018), .FEN(FEN[3884]), .op(N11018_t0) );
fim FAN_N11018_1 ( .fault(fault), .net(N11018), .FEN(FEN[3885]), .op(N11018_t1) );
fim FAN_N11056_0 ( .fault(fault), .net(N11056), .FEN(FEN[3886]), .op(N11056_t0) );
fim FAN_N11056_1 ( .fault(fault), .net(N11056), .FEN(FEN[3887]), .op(N11056_t1) );
fim FAN_N11059_0 ( .fault(fault), .net(N11059), .FEN(FEN[3888]), .op(N11059_t0) );
fim FAN_N11059_1 ( .fault(fault), .net(N11059), .FEN(FEN[3889]), .op(N11059_t1) );
fim FAN_N11067_0 ( .fault(fault), .net(N11067), .FEN(FEN[3890]), .op(N11067_t0) );
fim FAN_N11067_1 ( .fault(fault), .net(N11067), .FEN(FEN[3891]), .op(N11067_t1) );
fim FAN_N11070_0 ( .fault(fault), .net(N11070), .FEN(FEN[3892]), .op(N11070_t0) );
fim FAN_N11070_1 ( .fault(fault), .net(N11070), .FEN(FEN[3893]), .op(N11070_t1) );
fim FAN_N11044_0 ( .fault(fault), .net(N11044), .FEN(FEN[3894]), .op(N11044_t0) );
fim FAN_N11044_1 ( .fault(fault), .net(N11044), .FEN(FEN[3895]), .op(N11044_t1) );
fim FAN_N11047_0 ( .fault(fault), .net(N11047), .FEN(FEN[3896]), .op(N11047_t0) );
fim FAN_N11047_1 ( .fault(fault), .net(N11047), .FEN(FEN[3897]), .op(N11047_t1) );
fim FAN_N11050_0 ( .fault(fault), .net(N11050), .FEN(FEN[3898]), .op(N11050_t0) );
fim FAN_N11050_1 ( .fault(fault), .net(N11050), .FEN(FEN[3899]), .op(N11050_t1) );
fim FAN_N11053_0 ( .fault(fault), .net(N11053), .FEN(FEN[3900]), .op(N11053_t0) );
fim FAN_N11053_1 ( .fault(fault), .net(N11053), .FEN(FEN[3901]), .op(N11053_t1) );
fim FAN_N11062_0 ( .fault(fault), .net(N11062), .FEN(FEN[3902]), .op(N11062_t0) );
fim FAN_N11062_1 ( .fault(fault), .net(N11062), .FEN(FEN[3903]), .op(N11062_t1) );
fim FAN_N11103_0 ( .fault(fault), .net(N11103), .FEN(FEN[3904]), .op(N11103_t0) );
fim FAN_N11103_1 ( .fault(fault), .net(N11103), .FEN(FEN[3905]), .op(N11103_t1) );
fim FAN_N10283_0 ( .fault(fault), .net(N10283), .FEN(FEN[3906]), .op(N10283_t0) );
fim FAN_N10283_1 ( .fault(fault), .net(N10283), .FEN(FEN[3907]), .op(N10283_t1) );
fim FAN_N10283_2 ( .fault(fault), .net(N10283), .FEN(FEN[3908]), .op(N10283_t2) );
fim FAN_N11100_0 ( .fault(fault), .net(N11100), .FEN(FEN[3909]), .op(N11100_t0) );
fim FAN_N11100_1 ( .fault(fault), .net(N11100), .FEN(FEN[3910]), .op(N11100_t1) );
fim FAN_N11124_0 ( .fault(fault), .net(N11124), .FEN(FEN[3911]), .op(N11124_t0) );
fim FAN_N11124_1 ( .fault(fault), .net(N11124), .FEN(FEN[3912]), .op(N11124_t1) );
fim FAN_N11127_0 ( .fault(fault), .net(N11127), .FEN(FEN[3913]), .op(N11127_t0) );
fim FAN_N11127_1 ( .fault(fault), .net(N11127), .FEN(FEN[3914]), .op(N11127_t1) );
fim FAN_N11130_0 ( .fault(fault), .net(N11130), .FEN(FEN[3915]), .op(N11130_t0) );
fim FAN_N11130_1 ( .fault(fault), .net(N11130), .FEN(FEN[3916]), .op(N11130_t1) );
fim FAN_N11168_0 ( .fault(fault), .net(N11168), .FEN(FEN[3917]), .op(N11168_t0) );
fim FAN_N11168_1 ( .fault(fault), .net(N11168), .FEN(FEN[3918]), .op(N11168_t1) );
fim FAN_N11171_0 ( .fault(fault), .net(N11171), .FEN(FEN[3919]), .op(N11171_t0) );
fim FAN_N11171_1 ( .fault(fault), .net(N11171), .FEN(FEN[3920]), .op(N11171_t1) );
fim FAN_N11174_0 ( .fault(fault), .net(N11174), .FEN(FEN[3921]), .op(N11174_t0) );
fim FAN_N11174_1 ( .fault(fault), .net(N11174), .FEN(FEN[3922]), .op(N11174_t1) );
fim FAN_N11177_0 ( .fault(fault), .net(N11177), .FEN(FEN[3923]), .op(N11177_t0) );
fim FAN_N11177_1 ( .fault(fault), .net(N11177), .FEN(FEN[3924]), .op(N11177_t1) );
fim FAN_N11159_0 ( .fault(fault), .net(N11159), .FEN(FEN[3925]), .op(N11159_t0) );
fim FAN_N11159_1 ( .fault(fault), .net(N11159), .FEN(FEN[3926]), .op(N11159_t1) );
fim FAN_N1218_0 ( .fault(fault), .net(N1218), .FEN(FEN[3927]), .op(N1218_t0) );
fim FAN_N1218_1 ( .fault(fault), .net(N1218), .FEN(FEN[3928]), .op(N1218_t1) );
fim FAN_N1218_2 ( .fault(fault), .net(N1218), .FEN(FEN[3929]), .op(N1218_t2) );
fim FAN_N11156_0 ( .fault(fault), .net(N11156), .FEN(FEN[3930]), .op(N11156_t0) );
fim FAN_N11156_1 ( .fault(fault), .net(N11156), .FEN(FEN[3931]), .op(N11156_t1) );
fim FAN_N11165_0 ( .fault(fault), .net(N11165), .FEN(FEN[3932]), .op(N11165_t0) );
fim FAN_N11165_1 ( .fault(fault), .net(N11165), .FEN(FEN[3933]), .op(N11165_t1) );
fim FAN_N10497_0 ( .fault(fault), .net(N10497), .FEN(FEN[3934]), .op(N10497_t0) );
fim FAN_N10497_1 ( .fault(fault), .net(N10497), .FEN(FEN[3935]), .op(N10497_t1) );
fim FAN_N10497_2 ( .fault(fault), .net(N10497), .FEN(FEN[3936]), .op(N10497_t2) );
fim FAN_N11162_0 ( .fault(fault), .net(N11162), .FEN(FEN[3937]), .op(N11162_t0) );
fim FAN_N11162_1 ( .fault(fault), .net(N11162), .FEN(FEN[3938]), .op(N11162_t1) );
fim FAN_N11180_0 ( .fault(fault), .net(N11180), .FEN(FEN[3939]), .op(N11180_t0) );
fim FAN_N11180_1 ( .fault(fault), .net(N11180), .FEN(FEN[3940]), .op(N11180_t1) );
fim FAN_N11205_0 ( .fault(fault), .net(N11205), .FEN(FEN[3941]), .op(N11205_t0) );
fim FAN_N11205_1 ( .fault(fault), .net(N11205), .FEN(FEN[3942]), .op(N11205_t1) );
fim FAN_N11233_0 ( .fault(fault), .net(N11233), .FEN(FEN[3943]), .op(N11233_t0) );
fim FAN_N11233_1 ( .fault(fault), .net(N11233), .FEN(FEN[3944]), .op(N11233_t1) );
fim FAN_N11236_0 ( .fault(fault), .net(N11236), .FEN(FEN[3945]), .op(N11236_t0) );
fim FAN_N11236_1 ( .fault(fault), .net(N11236), .FEN(FEN[3946]), .op(N11236_t1) );
fim FAN_N11239_0 ( .fault(fault), .net(N11239), .FEN(FEN[3947]), .op(N11239_t0) );
fim FAN_N11239_1 ( .fault(fault), .net(N11239), .FEN(FEN[3948]), .op(N11239_t1) );
fim FAN_N11252_0 ( .fault(fault), .net(N11252), .FEN(FEN[3949]), .op(N11252_t0) );
fim FAN_N11252_1 ( .fault(fault), .net(N11252), .FEN(FEN[3950]), .op(N11252_t1) );
fim FAN_N11257_0 ( .fault(fault), .net(N11257), .FEN(FEN[3951]), .op(N11257_t0) );
fim FAN_N11257_1 ( .fault(fault), .net(N11257), .FEN(FEN[3952]), .op(N11257_t1) );
fim FAN_N11272_0 ( .fault(fault), .net(N11272), .FEN(FEN[3953]), .op(N11272_t0) );
fim FAN_N11272_1 ( .fault(fault), .net(N11272), .FEN(FEN[3954]), .op(N11272_t1) );
fim FAN_N11302_0 ( .fault(fault), .net(N11302), .FEN(FEN[3955]), .op(N11302_t0) );
fim FAN_N11302_1 ( .fault(fault), .net(N11302), .FEN(FEN[3956]), .op(N11302_t1) );
fim FAN_N11299_0 ( .fault(fault), .net(N11299), .FEN(FEN[3957]), .op(N11299_t0) );
fim FAN_N11299_1 ( .fault(fault), .net(N11299), .FEN(FEN[3958]), .op(N11299_t1) );
fim FAN_N11317_0 ( .fault(fault), .net(N11317), .FEN(FEN[3959]), .op(N11317_t0) );
fim FAN_N11317_1 ( .fault(fault), .net(N11317), .FEN(FEN[3960]), .op(N11317_t1) );
fim FAN_N11323_0 ( .fault(fault), .net(N11323), .FEN(FEN[3961]), .op(N11323_t0) );
fim FAN_N11323_1 ( .fault(fault), .net(N11323), .FEN(FEN[3962]), .op(N11323_t1) );
initial begin
    FEN <= {3962'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {3962'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,3962'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,3962'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN <= {FEN[3961:0], FEN[3962]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
// EndFaultModel

//Anchor
buf BUFF1_1 (N387, N1_t0);
buf BUFF1_2 (N388, N1_t1);
not NOT1_3 (N467, N57_t);
and AND2_4 (N469, N134_t, N133_t);
buf BUFF1_5 (N478, N248_t0);
buf BUFF1_6 (N482, N254_t0);
buf BUFF1_7 (N484, N257_t0);
buf BUFF1_8 (N486, N260_t0);
buf BUFF1_9 (N489, N263_t0);
buf BUFF1_10 (N492, N267_t0);
and AND4_11 (N494, N162_t, N172_t, N188_t, N199_t);
buf BUFF1_12 (N501, N274_t0);
buf BUFF1_13 (N505, N280_t0);
buf BUFF1_14 (N507, N283_t0);
buf BUFF1_15 (N509, N286_t0);
buf BUFF1_16 (N511, N289_t0);
buf BUFF1_17 (N513, N293_t0);
buf BUFF1_18 (N515, N296_t0);
buf BUFF1_19 (N517, N299_t0);
buf BUFF1_20 (N519, N303_t0);
and AND4_21 (N528, N150_t, N184_t, N228_t, N240_t);
buf BUFF1_22 (N535, N307_t0);
buf BUFF1_23 (N537, N310_t0);
buf BUFF1_24 (N539, N313_t0);
buf BUFF1_25 (N541, N316_t0);
buf BUFF1_26 (N543, N319_t0);
buf BUFF1_27 (N545, N322_t0);
buf BUFF1_28 (N547, N325_t0);
buf BUFF1_29 (N549, N328_t0);
buf BUFF1_30 (N551, N331_t0);
buf BUFF1_31 (N553, N334_t0);
buf BUFF1_32 (N556, N337_t0);
buf BUFF1_33 (N559, N343_t0);
buf BUFF1_34 (N561, N346_t0);
buf BUFF1_35 (N563, N349_t0);
buf BUFF1_36 (N565, N352_t0);
buf BUFF1_37 (N567, N355_t0);
buf BUFF1_38 (N569, N358_t0);
buf BUFF1_39 (N571, N361_t0);
buf BUFF1_40 (N573, N364_t0);
and AND4_41 (N575, N183_t, N182_t, N185_t, N186_t);
and AND4_42 (N578, N210_t, N152_t, N218_t, N230_t);
not NOT1_43 (N582, N15_t0);
not NOT1_44 (N585, N5_t0);
buf BUFF1_45 (N590, N1_t2);
not NOT1_46 (N593, N5_t1);
not NOT1_47 (N596, N5_t2);
not NOT1_48 (N599, N289_t1);
not NOT1_49 (N604, N299_t1);
not NOT1_50 (N609, N303_t1);
buf BUFF1_51 (N614, N38_t0);
buf BUFF1_52 (N625, N15_t1);
nand NAND2_53 (N628, N12_t0, N9_t0);
nand NAND2_54 (N632, N12_t1, N9_t1);
buf BUFF1_55 (N636, N38_t1);
not NOT1_56 (N641, N245_t0);
not NOT1_57 (N642, N248_t1);
buf BUFF1_58 (N643, N251_t0);
not NOT1_59 (N644, N251_t1);
not NOT1_60 (N651, N254_t1);
buf BUFF1_61 (N657, N106_t0);
not NOT1_62 (N660, N257_t1);
not NOT1_63 (N666, N260_t1);
not NOT1_64 (N672, N263_t1);
not NOT1_65 (N673, N267_t1);
not NOT1_66 (N674, N106_t1);
buf BUFF1_67 (N676, N18_t0);
buf BUFF1_68 (N682, N18_t1);
and AND2_69 (N688, N382_t0, N263_t2);
buf BUFF1_70 (N689, N18_t2);
not NOT1_71 (N695, N18_t3);
nand NAND2_72 (N700, N382_t1, N267_t2);
not NOT1_73 (N705, N271_t0);
not NOT1_74 (N706, N274_t1);
buf BUFF1_75 (N707, N277_t0);
not NOT1_76 (N708, N277_t1);
not NOT1_77 (N715, N280_t1);
not NOT1_78 (N721, N283_t1);
not NOT1_79 (N727, N286_t1);
not NOT1_80 (N733, N289_t2);
not NOT1_81 (N734, N293_t1);
not NOT1_82 (N742, N296_t1);
not NOT1_83 (N748, N299_t2);
not NOT1_84 (N749, N303_t2);
buf BUFF1_85 (N750, N367_t0);
not NOT1_86 (N758, N307_t1);
not NOT1_87 (N759, N310_t1);
not NOT1_88 (N762, N313_t1);
not NOT1_89 (N768, N316_t1);
not NOT1_90 (N774, N319_t1);
not NOT1_91 (N780, N322_t1);
not NOT1_92 (N786, N325_t1);
not NOT1_93 (N794, N328_t1);
not NOT1_94 (N800, N331_t1);
not NOT1_95 (N806, N334_t1);
not NOT1_96 (N812, N337_t1);
buf BUFF1_97 (N813, N340_t0);
not NOT1_98 (N814, N340_t1);
not NOT1_99 (N821, N343_t1);
not NOT1_100 (N827, N346_t1);
not NOT1_101 (N833, N349_t1);
not NOT1_102 (N839, N352_t1);
not NOT1_103 (N845, N355_t1);
not NOT1_104 (N853, N358_t1);
not NOT1_105 (N859, N361_t1);
not NOT1_106 (N865, N364_t1);
buf BUFF1_107 (N871, N367_t1);
nand NAND2_108 (N881, N467, N585);
not NOT1_109 (N882, N528_t0);
not NOT1_110 (N883, N578_t0);
not NOT1_111 (N884, N575_t0);
not NOT1_112 (N885, N494_t0);
and AND2_113 (N886, N528_t1, N578_t1);
and AND2_114 (N887, N575_t1, N494_t1);
buf BUFF1_115 (N889, N590_t0);
buf BUFF1_116 (N945, N657_t0);
not NOT1_117 (N957, N688);
and AND2_118 (N1028, N382_t2, N641);
nand NAND2_119 (N1029, N382_t3, N705);
and AND2_120 (N1109, N469_t0, N596_t0);
nand NAND2_121 (N1110, N242_t0, N593_t0);
not NOT1_122 (N1111, N625_t0);
nand NAND2_123 (N1112, N242_t1, N593_t1);
nand NAND2_124 (N1113, N469_t1, N596_t1);
not NOT1_125 (N1114, N625_t1);
not NOT1_126 (N1115, N871_t0);
buf BUFF1_127 (N1116, N590_t1);
buf BUFF1_128 (N1119, N628_t0);
buf BUFF1_129 (N1125, N682_t0);
buf BUFF1_130 (N1132, N628_t1);
buf BUFF1_131 (N1136, N682_t1);
buf BUFF1_132 (N1141, N628_t2);
buf BUFF1_133 (N1147, N682_t2);
buf BUFF1_134 (N1154, N632_t0);
buf BUFF1_135 (N1160, N676_t0);
and AND2_136 (N1167, N700_t0, N614_t0);
and AND2_137 (N1174, N700_t1, N614_t1);
buf BUFF1_138 (N1175, N682_t3);
buf BUFF1_139 (N1182, N676_t1);
not NOT1_140 (N1189, N657_t1);
not NOT1_141 (N1194, N676_t2);
not NOT1_142 (N1199, N682_t4);
not NOT1_143 (N1206, N689_t0);
buf BUFF1_144 (N1211, N695_t0);
not NOT1_145 (N1218, N750_t0);
not NOT1_146 (N1222, N1028);
buf BUFF1_147 (N1227, N632_t1);
buf BUFF1_148 (N1233, N676_t3);
buf BUFF1_149 (N1240, N632_t2);
buf BUFF1_150 (N1244, N676_t4);
buf BUFF1_151 (N1249, N689_t1);
buf BUFF1_152 (N1256, N689_t2);
buf BUFF1_153 (N1263, N695_t1);
buf BUFF1_154 (N1270, N689_t3);
buf BUFF1_155 (N1277, N689_t4);
buf BUFF1_156 (N1284, N700_t2);
buf BUFF1_157 (N1287, N614_t2);
buf BUFF1_158 (N1290, N666_t0);
buf BUFF1_159 (N1293, N660_t0);
buf BUFF1_160 (N1296, N651_t0);
buf BUFF1_161 (N1299, N614_t3);
buf BUFF1_162 (N1302, N644_t0);
buf BUFF1_163 (N1305, N700_t3);
buf BUFF1_164 (N1308, N614_t4);
buf BUFF1_165 (N1311, N614_t5);
buf BUFF1_166 (N1314, N666_t1);
buf BUFF1_167 (N1317, N660_t1);
buf BUFF1_168 (N1320, N651_t1);
buf BUFF1_169 (N1323, N644_t1);
buf BUFF1_170 (N1326, N609_t0);
buf BUFF1_171 (N1329, N604_t0);
buf BUFF1_172 (N1332, N742_t0);
buf BUFF1_173 (N1335, N599_t0);
buf BUFF1_174 (N1338, N727_t0);
buf BUFF1_175 (N1341, N721_t0);
buf BUFF1_176 (N1344, N715_t0);
buf BUFF1_177 (N1347, N734_t0);
buf BUFF1_178 (N1350, N708_t0);
buf BUFF1_179 (N1353, N609_t1);
buf BUFF1_180 (N1356, N604_t1);
buf BUFF1_181 (N1359, N742_t1);
buf BUFF1_182 (N1362, N734_t1);
buf BUFF1_183 (N1365, N599_t1);
buf BUFF1_184 (N1368, N727_t1);
buf BUFF1_185 (N1371, N721_t1);
buf BUFF1_186 (N1374, N715_t1);
buf BUFF1_187 (N1377, N708_t1);
buf BUFF1_188 (N1380, N806_t0);
buf BUFF1_189 (N1383, N800_t0);
buf BUFF1_190 (N1386, N794_t0);
buf BUFF1_191 (N1389, N786_t0);
buf BUFF1_192 (N1392, N780_t0);
buf BUFF1_193 (N1395, N774_t0);
buf BUFF1_194 (N1398, N768_t0);
buf BUFF1_195 (N1401, N762_t0);
buf BUFF1_196 (N1404, N806_t1);
buf BUFF1_197 (N1407, N800_t1);
buf BUFF1_198 (N1410, N794_t1);
buf BUFF1_199 (N1413, N780_t1);
buf BUFF1_200 (N1416, N774_t1);
buf BUFF1_201 (N1419, N768_t1);
buf BUFF1_202 (N1422, N762_t1);
buf BUFF1_203 (N1425, N786_t1);
buf BUFF1_204 (N1428, N636_t0);
buf BUFF1_205 (N1431, N636_t1);
buf BUFF1_206 (N1434, N865_t0);
buf BUFF1_207 (N1437, N859_t0);
buf BUFF1_208 (N1440, N853_t0);
buf BUFF1_209 (N1443, N845_t0);
buf BUFF1_210 (N1446, N839_t0);
buf BUFF1_211 (N1449, N833_t0);
buf BUFF1_212 (N1452, N827_t0);
buf BUFF1_213 (N1455, N821_t0);
buf BUFF1_214 (N1458, N814_t0);
buf BUFF1_215 (N1461, N865_t1);
buf BUFF1_216 (N1464, N859_t1);
buf BUFF1_217 (N1467, N853_t1);
buf BUFF1_218 (N1470, N839_t1);
buf BUFF1_219 (N1473, N833_t1);
buf BUFF1_220 (N1476, N827_t1);
buf BUFF1_221 (N1479, N821_t1);
buf BUFF1_222 (N1482, N845_t1);
buf BUFF1_223 (N1485, N814_t1);
not NOT1_224 (N1489, N1109);
buf BUFF1_225 (N1490, N1116_t0);
and AND2_226 (N1537, N957_t0, N614_t6);
and AND2_227 (N1551, N614_t7, N957_t1);
and AND2_228 (N1649, N1029_t0, N636_t2);
buf BUFF1_229 (N1703, N957_t2);
nor NOR2_230 (N1708, N957_t3, N614_t8);
buf BUFF1_231 (N1713, N957_t4);
nor NOR2_232 (N1721, N614_t9, N957_t5);
buf BUFF1_233 (N1758, N1029_t1);
and AND2_234 (N1781, N163_t, N1116_t1);
and AND2_235 (N1782, N170_t, N1125_t0);
not NOT1_236 (N1783, N1125_t1);
not NOT1_237 (N1789, N1136_t0);
and AND2_238 (N1793, N169_t, N1125_t2);
and AND2_239 (N1794, N168_t, N1125_t3);
and AND2_240 (N1795, N167_t, N1125_t4);
and AND2_241 (N1796, N166_t, N1136_t1);
and AND2_242 (N1797, N165_t, N1136_t2);
and AND2_243 (N1798, N164_t, N1136_t3);
not NOT1_244 (N1799, N1147_t0);
not NOT1_245 (N1805, N1160_t0);
and AND2_246 (N1811, N177_t, N1147_t1);
and AND2_247 (N1812, N176_t, N1147_t2);
and AND2_248 (N1813, N175_t, N1147_t3);
and AND2_249 (N1814, N174_t, N1147_t4);
and AND2_250 (N1815, N173_t, N1147_t5);
and AND2_251 (N1816, N157_t, N1160_t1);
and AND2_252 (N1817, N156_t, N1160_t2);
and AND2_253 (N1818, N155_t, N1160_t3);
and AND2_254 (N1819, N154_t, N1160_t4);
and AND2_255 (N1820, N153_t, N1160_t5);
not NOT1_256 (N1821, N1284_t0);
not NOT1_257 (N1822, N1287_t0);
not NOT1_258 (N1828, N1290_t0);
not NOT1_259 (N1829, N1293_t0);
not NOT1_260 (N1830, N1296_t0);
not NOT1_261 (N1832, N1299_t0);
not NOT1_262 (N1833, N1302_t0);
not NOT1_263 (N1834, N1305_t0);
not NOT1_264 (N1835, N1308_t0);
not NOT1_265 (N1839, N1311_t0);
not NOT1_266 (N1840, N1314_t0);
not NOT1_267 (N1841, N1317_t0);
not NOT1_268 (N1842, N1320_t0);
not NOT1_269 (N1843, N1323_t0);
not NOT1_270 (N1845, N1175_t0);
not NOT1_271 (N1851, N1182_t0);
and AND2_272 (N1857, N181_t, N1175_t1);
and AND2_273 (N1858, N171_t, N1175_t2);
and AND2_274 (N1859, N180_t, N1175_t3);
and AND2_275 (N1860, N179_t, N1175_t4);
and AND2_276 (N1861, N178_t, N1175_t5);
and AND2_277 (N1862, N161_t, N1182_t1);
and AND2_278 (N1863, N151_t, N1182_t2);
and AND2_279 (N1864, N160_t, N1182_t3);
and AND2_280 (N1865, N159_t, N1182_t4);
and AND2_281 (N1866, N158_t, N1182_t5);
not NOT1_282 (N1867, N1326_t0);
not NOT1_283 (N1868, N1329_t0);
not NOT1_284 (N1869, N1332_t0);
not NOT1_285 (N1870, N1335_t0);
not NOT1_286 (N1871, N1338_t0);
not NOT1_287 (N1872, N1341_t0);
not NOT1_288 (N1873, N1344_t0);
not NOT1_289 (N1874, N1347_t0);
not NOT1_290 (N1875, N1350_t0);
not NOT1_291 (N1876, N1353_t0);
not NOT1_292 (N1877, N1356_t0);
not NOT1_293 (N1878, N1359_t0);
not NOT1_294 (N1879, N1362_t0);
not NOT1_295 (N1880, N1365_t0);
not NOT1_296 (N1881, N1368_t0);
not NOT1_297 (N1882, N1371_t0);
not NOT1_298 (N1883, N1374_t0);
not NOT1_299 (N1884, N1377_t0);
buf BUFF1_300 (N1885, N1199_t0);
buf BUFF1_301 (N1892, N1194_t0);
buf BUFF1_302 (N1899, N1199_t1);
buf BUFF1_303 (N1906, N1194_t1);
not NOT1_304 (N1913, N1211_t0);
buf BUFF1_305 (N1919, N1194_t2);
and AND2_306 (N1926, N44_t0, N1211_t1);
and AND2_307 (N1927, N41_t0, N1211_t2);
and AND2_308 (N1928, N29_t0, N1211_t3);
and AND2_309 (N1929, N26_t0, N1211_t4);
and AND2_310 (N1930, N23_t0, N1211_t5);
not NOT1_311 (N1931, N1380_t0);
not NOT1_312 (N1932, N1383_t0);
not NOT1_313 (N1933, N1386_t0);
not NOT1_314 (N1934, N1389_t0);
not NOT1_315 (N1935, N1392_t0);
not NOT1_316 (N1936, N1395_t0);
not NOT1_317 (N1937, N1398_t0);
not NOT1_318 (N1938, N1401_t0);
not NOT1_319 (N1939, N1404_t0);
not NOT1_320 (N1940, N1407_t0);
not NOT1_321 (N1941, N1410_t0);
not NOT1_322 (N1942, N1413_t0);
not NOT1_323 (N1943, N1416_t0);
not NOT1_324 (N1944, N1419_t0);
not NOT1_325 (N1945, N1422_t0);
not NOT1_326 (N1946, N1425_t0);
not NOT1_327 (N1947, N1233_t0);
not NOT1_328 (N1953, N1244_t0);
and AND2_329 (N1957, N209_t, N1233_t1);
and AND2_330 (N1958, N216_t, N1233_t2);
and AND2_331 (N1959, N215_t, N1233_t3);
and AND2_332 (N1960, N214_t, N1233_t4);
and AND2_333 (N1961, N213_t, N1244_t1);
and AND2_334 (N1962, N212_t, N1244_t2);
and AND2_335 (N1963, N211_t, N1244_t3);
not NOT1_336 (N1965, N1428_t0);
and AND2_337 (N1966, N1222_t0, N636_t3);
not NOT1_338 (N1967, N1431_t0);
not NOT1_339 (N1968, N1434_t0);
not NOT1_340 (N1969, N1437_t0);
not NOT1_341 (N1970, N1440_t0);
not NOT1_342 (N1971, N1443_t0);
not NOT1_343 (N1972, N1446_t0);
not NOT1_344 (N1973, N1449_t0);
not NOT1_345 (N1974, N1452_t0);
not NOT1_346 (N1975, N1455_t0);
not NOT1_347 (N1976, N1458_t0);
not NOT1_348 (N1977, N1249_t0);
not NOT1_349 (N1983, N1256_t0);
and AND2_350 (N1989, N642, N1249_t1);
and AND2_351 (N1990, N644_t2, N1249_t2);
and AND2_352 (N1991, N651_t2, N1249_t3);
and AND2_353 (N1992, N674, N1249_t4);
and AND2_354 (N1993, N660_t2, N1249_t5);
and AND2_355 (N1994, N666_t2, N1256_t1);
and AND2_356 (N1995, N672, N1256_t2);
and AND2_357 (N1996, N673, N1256_t3);
not NOT1_358 (N1997, N1263_t0);
buf BUFF1_359 (N2003, N1194_t3);
and AND2_360 (N2010, N47_t0, N1263_t1);
and AND2_361 (N2011, N35_t0, N1263_t2);
and AND2_362 (N2012, N32_t0, N1263_t3);
and AND2_363 (N2013, N50_t0, N1263_t4);
and AND2_364 (N2014, N66_t0, N1263_t5);
not NOT1_365 (N2015, N1461_t0);
not NOT1_366 (N2016, N1464_t0);
not NOT1_367 (N2017, N1467_t0);
not NOT1_368 (N2018, N1470_t0);
not NOT1_369 (N2019, N1473_t0);
not NOT1_370 (N2020, N1476_t0);
not NOT1_371 (N2021, N1479_t0);
not NOT1_372 (N2022, N1482_t0);
not NOT1_373 (N2023, N1485_t0);
buf BUFF1_374 (N2024, N1206_t0);
buf BUFF1_375 (N2031, N1206_t1);
buf BUFF1_376 (N2038, N1206_t2);
buf BUFF1_377 (N2045, N1206_t3);
not NOT1_378 (N2052, N1270_t0);
not NOT1_379 (N2058, N1277_t0);
and AND2_380 (N2064, N706, N1270_t1);
and AND2_381 (N2065, N708_t2, N1270_t2);
and AND2_382 (N2066, N715_t2, N1270_t3);
and AND2_383 (N2067, N721_t2, N1270_t4);
and AND2_384 (N2068, N727_t2, N1270_t5);
and AND2_385 (N2069, N733, N1277_t1);
and AND2_386 (N2070, N734_t2, N1277_t2);
and AND2_387 (N2071, N742_t2, N1277_t3);
and AND2_388 (N2072, N748, N1277_t4);
and AND2_389 (N2073, N749, N1277_t5);
buf BUFF1_390 (N2074, N1189_t0);
buf BUFF1_391 (N2081, N1189_t1);
buf BUFF1_392 (N2086, N1222_t1);
nand NAND2_393 (N2107, N1287_t1, N1821);
nand NAND2_394 (N2108, N1284_t1, N1822);
not NOT1_395 (N2110, N1703_t0);
nand NAND2_396 (N2111, N1703_t1, N1832);
nand NAND2_397 (N2112, N1308_t1, N1834);
nand NAND2_398 (N2113, N1305_t1, N1835);
not NOT1_399 (N2114, N1713_t0);
nand NAND2_400 (N2115, N1713_t1, N1839);
not NOT1_401 (N2117, N1721_t0);
not NOT1_402 (N2171, N1758_t0);
nand NAND2_403 (N2172, N1758_t1, N1965);
not NOT1_404 (N2230, N1708_t0);
buf BUFF1_405 (N2231, N1537_t0);
buf BUFF1_406 (N2235, N1551_t0);
or OR2_407 (N2239, N1783_t0, N1782);
or OR2_408 (N2240, N1783_t1, N1125_t5);
or OR2_409 (N2241, N1783_t2, N1793);
or OR2_410 (N2242, N1783_t3, N1794);
or OR2_411 (N2243, N1783_t4, N1795);
or OR2_412 (N2244, N1789_t0, N1796);
or OR2_413 (N2245, N1789_t1, N1797);
or OR2_414 (N2246, N1789_t2, N1798);
or OR2_415 (N2247, N1799_t0, N1811);
or OR2_416 (N2248, N1799_t1, N1812);
or OR2_417 (N2249, N1799_t2, N1813);
or OR2_418 (N2250, N1799_t3, N1814);
or OR2_419 (N2251, N1799_t4, N1815);
or OR2_420 (N2252, N1805_t0, N1816);
or OR2_421 (N2253, N1805_t1, N1817);
or OR2_422 (N2254, N1805_t2, N1818);
or OR2_423 (N2255, N1805_t3, N1819);
or OR2_424 (N2256, N1805_t4, N1820);
nand NAND2_425 (N2257, N2107, N2108);
not NOT1_426 (N2267, N2074_t0);
nand NAND2_427 (N2268, N1299_t1, N2110);
nand NAND2_428 (N2269, N2112, N2113);
nand NAND2_429 (N2274, N1311_t1, N2114);
not NOT1_430 (N2275, N2081_t0);
and AND2_431 (N2277, N141_t0, N1845_t0);
and AND2_432 (N2278, N147_t0, N1845_t1);
and AND2_433 (N2279, N138_t0, N1845_t2);
and AND2_434 (N2280, N144_t0, N1845_t3);
and AND2_435 (N2281, N135_t0, N1845_t4);
and AND2_436 (N2282, N141_t1, N1851_t0);
and AND2_437 (N2283, N147_t1, N1851_t1);
and AND2_438 (N2284, N138_t1, N1851_t2);
and AND2_439 (N2285, N144_t1, N1851_t3);
and AND2_440 (N2286, N135_t1, N1851_t4);
not NOT1_441 (N2287, N1885_t0);
not NOT1_442 (N2293, N1892_t0);
and AND2_443 (N2299, N103_t0, N1885_t1);
and AND2_444 (N2300, N130_t0, N1885_t2);
and AND2_445 (N2301, N127_t0, N1885_t3);
and AND2_446 (N2302, N124_t0, N1885_t4);
and AND2_447 (N2303, N100_t0, N1885_t5);
and AND2_448 (N2304, N103_t1, N1892_t1);
and AND2_449 (N2305, N130_t1, N1892_t2);
and AND2_450 (N2306, N127_t1, N1892_t3);
and AND2_451 (N2307, N124_t1, N1892_t4);
and AND2_452 (N2308, N100_t1, N1892_t5);
not NOT1_453 (N2309, N1899_t0);
not NOT1_454 (N2315, N1906_t0);
and AND2_455 (N2321, N115_t0, N1899_t1);
and AND2_456 (N2322, N118_t0, N1899_t2);
and AND2_457 (N2323, N97_t0, N1899_t3);
and AND2_458 (N2324, N94_t0, N1899_t4);
and AND2_459 (N2325, N121_t0, N1899_t5);
and AND2_460 (N2326, N115_t1, N1906_t1);
and AND2_461 (N2327, N118_t1, N1906_t2);
and AND2_462 (N2328, N97_t1, N1906_t3);
and AND2_463 (N2329, N94_t1, N1906_t4);
and AND2_464 (N2330, N121_t1, N1906_t5);
not NOT1_465 (N2331, N1919_t0);
and AND2_466 (N2337, N208_t, N1913_t0);
and AND2_467 (N2338, N198_t, N1913_t1);
and AND2_468 (N2339, N207_t, N1913_t2);
and AND2_469 (N2340, N206_t, N1913_t3);
and AND2_470 (N2341, N205_t, N1913_t4);
and AND2_471 (N2342, N44_t1, N1919_t1);
and AND2_472 (N2343, N41_t1, N1919_t2);
and AND2_473 (N2344, N29_t1, N1919_t3);
and AND2_474 (N2345, N26_t1, N1919_t4);
and AND2_475 (N2346, N23_t1, N1919_t5);
or OR2_476 (N2347, N1947_t0, N1233_t5);
or OR2_477 (N2348, N1947_t1, N1957);
or OR2_478 (N2349, N1947_t2, N1958);
or OR2_479 (N2350, N1947_t3, N1959);
or OR2_480 (N2351, N1947_t4, N1960);
or OR2_481 (N2352, N1953_t0, N1961);
or OR2_482 (N2353, N1953_t1, N1962);
or OR2_483 (N2354, N1953_t2, N1963);
nand NAND2_484 (N2355, N1428_t1, N2171);
not NOT1_485 (N2356, N2086_t0);
nand NAND2_486 (N2357, N2086_t1, N1967);
and AND2_487 (N2358, N114_t, N1977_t0);
and AND2_488 (N2359, N113_t, N1977_t1);
and AND2_489 (N2360, N111_t, N1977_t2);
and AND2_490 (N2361, N87_t, N1977_t3);
and AND2_491 (N2362, N112_t, N1977_t4);
and AND2_492 (N2363, N88_t, N1983_t0);
and AND2_493 (N2364, N245_t1, N1983_t1);
and AND2_494 (N2365, N271_t1, N1983_t2);
and AND2_495 (N2366, N759_t0, N1983_t3);
and AND2_496 (N2367, N70_t0, N1983_t4);
not NOT1_497 (N2368, N2003_t0);
and AND2_498 (N2374, N193_t, N1997_t0);
and AND2_499 (N2375, N192_t, N1997_t1);
and AND2_500 (N2376, N191_t, N1997_t2);
and AND2_501 (N2377, N190_t, N1997_t3);
and AND2_502 (N2378, N189_t, N1997_t4);
and AND2_503 (N2379, N47_t1, N2003_t1);
and AND2_504 (N2380, N35_t1, N2003_t2);
and AND2_505 (N2381, N32_t1, N2003_t3);
and AND2_506 (N2382, N50_t1, N2003_t4);
and AND2_507 (N2383, N66_t1, N2003_t5);
not NOT1_508 (N2384, N2024_t0);
not NOT1_509 (N2390, N2031_t0);
and AND2_510 (N2396, N58_t, N2024_t1);
and AND2_511 (N2397, N77_t, N2024_t2);
and AND2_512 (N2398, N78_t, N2024_t3);
and AND2_513 (N2399, N59_t, N2024_t4);
and AND2_514 (N2400, N81_t, N2024_t5);
and AND2_515 (N2401, N80_t, N2031_t1);
and AND2_516 (N2402, N79_t, N2031_t2);
and AND2_517 (N2403, N60_t, N2031_t3);
and AND2_518 (N2404, N61_t, N2031_t4);
and AND2_519 (N2405, N62_t, N2031_t5);
not NOT1_520 (N2406, N2038_t0);
not NOT1_521 (N2412, N2045_t0);
and AND2_522 (N2418, N69_t, N2038_t1);
and AND2_523 (N2419, N70_t1, N2038_t2);
and AND2_524 (N2420, N74_t, N2038_t3);
and AND2_525 (N2421, N76_t, N2038_t4);
and AND2_526 (N2422, N75_t, N2038_t5);
and AND2_527 (N2423, N73_t, N2045_t1);
and AND2_528 (N2424, N53_t, N2045_t2);
and AND2_529 (N2425, N54_t, N2045_t3);
and AND2_530 (N2426, N55_t, N2045_t4);
and AND2_531 (N2427, N56_t, N2045_t5);
and AND2_532 (N2428, N82_t, N2052_t0);
and AND2_533 (N2429, N65_t, N2052_t1);
and AND2_534 (N2430, N83_t, N2052_t2);
and AND2_535 (N2431, N84_t, N2052_t3);
and AND2_536 (N2432, N85_t, N2052_t4);
and AND2_537 (N2433, N64_t, N2058_t0);
and AND2_538 (N2434, N63_t, N2058_t1);
and AND2_539 (N2435, N86_t, N2058_t2);
and AND2_540 (N2436, N109_t, N2058_t3);
and AND2_541 (N2437, N110_t, N2058_t4);
and AND2_542 (N2441, N2239, N1119_t0);
and AND2_543 (N2442, N2240, N1119_t1);
and AND2_544 (N2446, N2241, N1119_t2);
and AND2_545 (N2450, N2242, N1119_t3);
and AND2_546 (N2454, N2243, N1119_t4);
and AND2_547 (N2458, N2244, N1132_t0);
and AND2_548 (N2462, N2247, N1141_t0);
and AND2_549 (N2466, N2248, N1141_t1);
and AND2_550 (N2470, N2249, N1141_t2);
and AND2_551 (N2474, N2250, N1141_t3);
and AND2_552 (N2478, N2251, N1141_t4);
and AND2_553 (N2482, N2252, N1154_t0);
and AND2_554 (N2488, N2253, N1154_t1);
and AND2_555 (N2496, N2254, N1154_t2);
and AND2_556 (N2502, N2255, N1154_t3);
and AND2_557 (N2508, N2256, N1154_t4);
nand NAND2_558 (N2523, N2268, N2111);
nand NAND2_559 (N2533, N2274, N2115);
not NOT1_560 (N2537, N2235_t0);
or OR2_561 (N2538, N2278, N1858);
or OR2_562 (N2542, N2279, N1859);
or OR2_563 (N2546, N2280, N1860);
or OR2_564 (N2550, N2281, N1861);
or OR2_565 (N2554, N2283, N1863);
or OR2_566 (N2561, N2284, N1864);
or OR2_567 (N2567, N2285, N1865);
or OR2_568 (N2573, N2286, N1866);
or OR2_569 (N2604, N2338, N1927);
or OR2_570 (N2607, N2339, N1928);
or OR2_571 (N2611, N2340, N1929);
or OR2_572 (N2615, N2341, N1930);
and AND2_573 (N2619, N2348, N1227_t0);
and AND2_574 (N2626, N2349, N1227_t1);
and AND2_575 (N2632, N2350, N1227_t2);
and AND2_576 (N2638, N2351, N1227_t3);
and AND2_577 (N2644, N2352, N1240_t0);
nand NAND2_578 (N2650, N2355, N2172);
nand NAND2_579 (N2653, N1431_t1, N2356);
or OR2_580 (N2654, N2359, N1990);
or OR2_581 (N2658, N2360, N1991);
or OR2_582 (N2662, N2361, N1992);
or OR2_583 (N2666, N2362, N1993);
or OR2_584 (N2670, N2363, N1994);
or OR2_585 (N2674, N2366, N1256_t4);
or OR2_586 (N2680, N2367, N1256_t5);
or OR2_587 (N2688, N2374, N2010);
or OR2_588 (N2692, N2375, N2011);
or OR2_589 (N2696, N2376, N2012);
or OR2_590 (N2700, N2377, N2013);
or OR2_591 (N2704, N2378, N2014);
and AND2_592 (N2728, N2347, N1227_t4);
or OR2_593 (N2729, N2429, N2065);
or OR2_594 (N2733, N2430, N2066);
or OR2_595 (N2737, N2431, N2067);
or OR2_596 (N2741, N2432, N2068);
or OR2_597 (N2745, N2433, N2069);
or OR2_598 (N2749, N2434, N2070);
or OR2_599 (N2753, N2435, N2071);
or OR2_600 (N2757, N2436, N2072);
or OR2_601 (N2761, N2437, N2073);
not NOT1_602 (N2765, N2231_t0);
and AND2_603 (N2766, N2354, N1240_t1);
and AND2_604 (N2769, N2353, N1240_t2);
and AND2_605 (N2772, N2246, N1132_t1);
and AND2_606 (N2775, N2245, N1132_t2);
or OR2_607 (N2778, N2282, N1862);
or OR2_608 (N2781, N2358, N1989);
or OR2_609 (N2784, N2365, N1996);
or OR2_610 (N2787, N2364, N1995);
or OR2_611 (N2790, N2337, N1926);
or OR2_612 (N2793, N2277, N1857);
or OR2_613 (N2796, N2428, N2064);
and AND2_614 (N2866, N2257_t0, N1537_t1);
and AND2_615 (N2867, N2257_t1, N1537_t2);
and AND2_616 (N2868, N2257_t2, N1537_t3);
and AND2_617 (N2869, N2257_t3, N1537_t4);
and AND2_618 (N2878, N2269_t0, N1551_t1);
and AND2_619 (N2913, N204_t, N2287_t0);
and AND2_620 (N2914, N203_t, N2287_t1);
and AND2_621 (N2915, N202_t, N2287_t2);
and AND2_622 (N2916, N201_t, N2287_t3);
and AND2_623 (N2917, N200_t, N2287_t4);
and AND2_624 (N2918, N235_t, N2293_t0);
and AND2_625 (N2919, N234_t, N2293_t1);
and AND2_626 (N2920, N233_t, N2293_t2);
and AND2_627 (N2921, N232_t, N2293_t3);
and AND2_628 (N2922, N231_t, N2293_t4);
and AND2_629 (N2923, N197_t, N2309_t0);
and AND2_630 (N2924, N187_t, N2309_t1);
and AND2_631 (N2925, N196_t, N2309_t2);
and AND2_632 (N2926, N195_t, N2309_t3);
and AND2_633 (N2927, N194_t, N2309_t4);
and AND2_634 (N2928, N227_t, N2315_t0);
and AND2_635 (N2929, N217_t, N2315_t1);
and AND2_636 (N2930, N226_t, N2315_t2);
and AND2_637 (N2931, N225_t, N2315_t3);
and AND2_638 (N2932, N224_t, N2315_t4);
and AND2_639 (N2933, N239_t, N2331_t0);
and AND2_640 (N2934, N229_t, N2331_t1);
and AND2_641 (N2935, N238_t, N2331_t2);
and AND2_642 (N2936, N237_t, N2331_t3);
and AND2_643 (N2937, N236_t, N2331_t4);
nand NAND2_644 (N2988, N2653, N2357);
and AND2_645 (N3005, N223_t, N2368_t0);
and AND2_646 (N3006, N222_t, N2368_t1);
and AND2_647 (N3007, N221_t, N2368_t2);
and AND2_648 (N3008, N220_t, N2368_t3);
and AND2_649 (N3009, N219_t, N2368_t4);
and AND2_650 (N3020, N812, N2384_t0);
and AND2_651 (N3021, N814_t2, N2384_t1);
and AND2_652 (N3022, N821_t2, N2384_t2);
and AND2_653 (N3023, N827_t2, N2384_t3);
and AND2_654 (N3024, N833_t2, N2384_t4);
and AND2_655 (N3025, N839_t2, N2390_t0);
and AND2_656 (N3026, N845_t2, N2390_t1);
and AND2_657 (N3027, N853_t2, N2390_t2);
and AND2_658 (N3028, N859_t2, N2390_t3);
and AND2_659 (N3029, N865_t2, N2390_t4);
and AND2_660 (N3032, N758, N2406_t0);
and AND2_661 (N3033, N759_t1, N2406_t1);
and AND2_662 (N3034, N762_t2, N2406_t2);
and AND2_663 (N3035, N768_t2, N2406_t3);
and AND2_664 (N3036, N774_t2, N2406_t4);
and AND2_665 (N3037, N780_t2, N2412_t0);
and AND2_666 (N3038, N786_t2, N2412_t1);
and AND2_667 (N3039, N794_t2, N2412_t2);
and AND2_668 (N3040, N800_t2, N2412_t3);
and AND2_669 (N3041, N806_t2, N2412_t4);
buf BUFF1_670 (N3061, N2257_t4);
buf BUFF1_671 (N3064, N2257_t5);
buf BUFF1_672 (N3067, N2269_t1);
buf BUFF1_673 (N3070, N2269_t2);
not NOT1_674 (N3073, N2728);
not NOT1_675 (N3080, N2441);
and AND2_676 (N3096, N666_t3, N2644_t0);
and AND2_677 (N3097, N660_t3, N2638_t0);
and AND2_678 (N3101, N1189_t2, N2632_t0);
and AND2_679 (N3107, N651_t3, N2626_t0);
and AND2_680 (N3114, N644_t3, N2619_t0);
and AND2_681 (N3122, N2523_t0, N2257_t6);
or OR2_682 (N3126, N1167_t0, N2866);
and AND2_683 (N3130, N2523_t1, N2257_t7);
or OR2_684 (N3131, N1167_t1, N2869);
and AND2_685 (N3134, N2523_t2, N2257_t8);
not NOT1_686 (N3135, N2533_t0);
and AND2_687 (N3136, N666_t4, N2644_t1);
and AND2_688 (N3137, N660_t4, N2638_t1);
and AND2_689 (N3140, N1189_t3, N2632_t1);
and AND2_690 (N3144, N651_t4, N2626_t1);
and AND2_691 (N3149, N644_t4, N2619_t1);
and AND2_692 (N3155, N2533_t1, N2269_t3);
or OR2_693 (N3159, N1174, N2878);
not NOT1_694 (N3167, N2778_t0);
and AND2_695 (N3168, N609_t2, N2508_t0);
and AND2_696 (N3169, N604_t2, N2502_t0);
and AND2_697 (N3173, N742_t3, N2496_t0);
and AND2_698 (N3178, N734_t3, N2488_t0);
and AND2_699 (N3184, N599_t2, N2482_t0);
and AND2_700 (N3185, N727_t3, N2573_t0);
and AND2_701 (N3189, N721_t3, N2567_t0);
and AND2_702 (N3195, N715_t3, N2561_t0);
and AND2_703 (N3202, N708_t3, N2554_t0);
and AND2_704 (N3210, N609_t3, N2508_t1);
and AND2_705 (N3211, N604_t3, N2502_t1);
and AND2_706 (N3215, N742_t4, N2496_t1);
and AND2_707 (N3221, N2488_t1, N734_t4);
and AND2_708 (N3228, N599_t3, N2482_t1);
and AND2_709 (N3229, N727_t4, N2573_t1);
and AND2_710 (N3232, N721_t4, N2567_t1);
and AND2_711 (N3236, N715_t4, N2561_t1);
and AND2_712 (N3241, N708_t4, N2554_t1);
or OR2_713 (N3247, N2913, N2299);
or OR2_714 (N3251, N2914, N2300);
or OR2_715 (N3255, N2915, N2301);
or OR2_716 (N3259, N2916, N2302);
or OR2_717 (N3263, N2917, N2303);
or OR2_718 (N3267, N2918, N2304);
or OR2_719 (N3273, N2919, N2305);
or OR2_720 (N3281, N2920, N2306);
or OR2_721 (N3287, N2921, N2307);
or OR2_722 (N3293, N2922, N2308);
or OR2_723 (N3299, N2924, N2322);
or OR2_724 (N3303, N2925, N2323);
or OR2_725 (N3307, N2926, N2324);
or OR2_726 (N3311, N2927, N2325);
or OR2_727 (N3315, N2929, N2327);
or OR2_728 (N3322, N2930, N2328);
or OR2_729 (N3328, N2931, N2329);
or OR2_730 (N3334, N2932, N2330);
or OR2_731 (N3340, N2934, N2343);
or OR2_732 (N3343, N2935, N2344);
or OR2_733 (N3349, N2936, N2345);
or OR2_734 (N3355, N2937, N2346);
and AND2_735 (N3361, N2761_t0, N2478_t0);
and AND2_736 (N3362, N2757_t0, N2474_t0);
and AND2_737 (N3363, N2753_t0, N2470_t0);
and AND2_738 (N3364, N2749_t0, N2466_t0);
and AND2_739 (N3365, N2745_t0, N2462_t0);
and AND2_740 (N3366, N2741_t0, N2550_t0);
and AND2_741 (N3367, N2737_t0, N2546_t0);
and AND2_742 (N3368, N2733_t0, N2542_t0);
and AND2_743 (N3369, N2729_t0, N2538_t0);
and AND2_744 (N3370, N2670_t0, N2458_t0);
and AND2_745 (N3371, N2666_t0, N2454_t0);
and AND2_746 (N3372, N2662_t0, N2450_t0);
and AND2_747 (N3373, N2658_t0, N2446_t0);
and AND2_748 (N3374, N2654_t0, N2442_t0);
and AND2_749 (N3375, N2988, N2650_t0);
and AND2_750 (N3379, N2650_t1, N1966);
not NOT1_751 (N3380, N2781_t0);
and AND2_752 (N3381, N695_t2, N2604_t0);
or OR2_753 (N3384, N3005, N2379);
or OR2_754 (N3390, N3006, N2380);
or OR2_755 (N3398, N3007, N2381);
or OR2_756 (N3404, N3008, N2382);
or OR2_757 (N3410, N3009, N2383);
or OR2_758 (N3416, N3021, N2397);
or OR2_759 (N3420, N3022, N2398);
or OR2_760 (N3424, N3023, N2399);
or OR2_761 (N3428, N3024, N2400);
or OR2_762 (N3432, N3025, N2401);
or OR2_763 (N3436, N3026, N2402);
or OR2_764 (N3440, N3027, N2403);
or OR2_765 (N3444, N3028, N2404);
or OR2_766 (N3448, N3029, N2405);
not NOT1_767 (N3452, N2790_t0);
not NOT1_768 (N3453, N2793_t0);
or OR2_769 (N3454, N3034, N2420);
or OR2_770 (N3458, N3035, N2421);
or OR2_771 (N3462, N3036, N2422);
or OR2_772 (N3466, N3037, N2423);
or OR2_773 (N3470, N3038, N2424);
or OR2_774 (N3474, N3039, N2425);
or OR2_775 (N3478, N3040, N2426);
or OR2_776 (N3482, N3041, N2427);
not NOT1_777 (N3486, N2796_t0);
buf BUFF1_778 (N3487, N2644_t2);
buf BUFF1_779 (N3490, N2638_t2);
buf BUFF1_780 (N3493, N2632_t2);
buf BUFF1_781 (N3496, N2626_t2);
buf BUFF1_782 (N3499, N2619_t2);
buf BUFF1_783 (N3502, N2523_t3);
nor NOR2_784 (N3507, N1167_t2, N2868);
buf BUFF1_785 (N3510, N2523_t4);
nor NOR2_786 (N3515, N644_t5, N2619_t3);
buf BUFF1_787 (N3518, N2644_t3);
buf BUFF1_788 (N3521, N2638_t3);
buf BUFF1_789 (N3524, N2632_t3);
buf BUFF1_790 (N3527, N2626_t3);
buf BUFF1_791 (N3530, N2619_t4);
buf BUFF1_792 (N3535, N2619_t5);
buf BUFF1_793 (N3539, N2632_t4);
buf BUFF1_794 (N3542, N2626_t4);
buf BUFF1_795 (N3545, N2644_t4);
buf BUFF1_796 (N3548, N2638_t4);
not NOT1_797 (N3551, N2766_t0);
not NOT1_798 (N3552, N2769_t0);
buf BUFF1_799 (N3553, N2442_t1);
buf BUFF1_800 (N3557, N2450_t1);
buf BUFF1_801 (N3560, N2446_t1);
buf BUFF1_802 (N3563, N2458_t1);
buf BUFF1_803 (N3566, N2454_t1);
not NOT1_804 (N3569, N2772_t0);
not NOT1_805 (N3570, N2775_t0);
buf BUFF1_806 (N3571, N2554_t2);
buf BUFF1_807 (N3574, N2567_t2);
buf BUFF1_808 (N3577, N2561_t2);
buf BUFF1_809 (N3580, N2482_t2);
buf BUFF1_810 (N3583, N2573_t2);
buf BUFF1_811 (N3586, N2496_t2);
buf BUFF1_812 (N3589, N2488_t2);
buf BUFF1_813 (N3592, N2508_t2);
buf BUFF1_814 (N3595, N2502_t2);
buf BUFF1_815 (N3598, N2508_t3);
buf BUFF1_816 (N3601, N2502_t3);
buf BUFF1_817 (N3604, N2496_t3);
buf BUFF1_818 (N3607, N2482_t3);
buf BUFF1_819 (N3610, N2573_t3);
buf BUFF1_820 (N3613, N2567_t3);
buf BUFF1_821 (N3616, N2561_t3);
buf BUFF1_822 (N3619, N2488_t3);
buf BUFF1_823 (N3622, N2554_t3);
nor NOR2_824 (N3625, N734_t5, N2488_t4);
nor NOR2_825 (N3628, N708_t5, N2554_t4);
buf BUFF1_826 (N3631, N2508_t4);
buf BUFF1_827 (N3634, N2502_t4);
buf BUFF1_828 (N3637, N2496_t4);
buf BUFF1_829 (N3640, N2488_t5);
buf BUFF1_830 (N3643, N2482_t4);
buf BUFF1_831 (N3646, N2573_t4);
buf BUFF1_832 (N3649, N2567_t4);
buf BUFF1_833 (N3652, N2561_t4);
buf BUFF1_834 (N3655, N2554_t5);
nor NOR2_835 (N3658, N2488_t6, N734_t6);
buf BUFF1_836 (N3661, N2674_t0);
buf BUFF1_837 (N3664, N2674_t1);
buf BUFF1_838 (N3667, N2761_t1);
buf BUFF1_839 (N3670, N2478_t1);
buf BUFF1_840 (N3673, N2757_t1);
buf BUFF1_841 (N3676, N2474_t1);
buf BUFF1_842 (N3679, N2753_t1);
buf BUFF1_843 (N3682, N2470_t1);
buf BUFF1_844 (N3685, N2745_t1);
buf BUFF1_845 (N3688, N2462_t1);
buf BUFF1_846 (N3691, N2741_t1);
buf BUFF1_847 (N3694, N2550_t1);
buf BUFF1_848 (N3697, N2737_t1);
buf BUFF1_849 (N3700, N2546_t1);
buf BUFF1_850 (N3703, N2733_t1);
buf BUFF1_851 (N3706, N2542_t1);
buf BUFF1_852 (N3709, N2749_t1);
buf BUFF1_853 (N3712, N2466_t1);
buf BUFF1_854 (N3715, N2729_t1);
buf BUFF1_855 (N3718, N2538_t1);
buf BUFF1_856 (N3721, N2704_t0);
buf BUFF1_857 (N3724, N2700_t0);
buf BUFF1_858 (N3727, N2696_t0);
buf BUFF1_859 (N3730, N2688_t0);
buf BUFF1_860 (N3733, N2692_t0);
buf BUFF1_861 (N3736, N2670_t1);
buf BUFF1_862 (N3739, N2458_t2);
buf BUFF1_863 (N3742, N2666_t1);
buf BUFF1_864 (N3745, N2454_t2);
buf BUFF1_865 (N3748, N2662_t1);
buf BUFF1_866 (N3751, N2450_t2);
buf BUFF1_867 (N3754, N2658_t1);
buf BUFF1_868 (N3757, N2446_t2);
buf BUFF1_869 (N3760, N2654_t1);
buf BUFF1_870 (N3763, N2442_t2);
buf BUFF1_871 (N3766, N2654_t2);
buf BUFF1_872 (N3769, N2662_t2);
buf BUFF1_873 (N3772, N2658_t2);
buf BUFF1_874 (N3775, N2670_t2);
buf BUFF1_875 (N3778, N2666_t2);
not NOT1_876 (N3781, N2784_t0);
not NOT1_877 (N3782, N2787_t0);
or OR2_878 (N3783, N2928, N2326);
or OR2_879 (N3786, N2933, N2342);
or OR2_880 (N3789, N2923, N2321);
buf BUFF1_881 (N3792, N2688_t1);
buf BUFF1_882 (N3795, N2696_t1);
buf BUFF1_883 (N3798, N2692_t1);
buf BUFF1_884 (N3801, N2704_t1);
buf BUFF1_885 (N3804, N2700_t1);
buf BUFF1_886 (N3807, N2604_t1);
buf BUFF1_887 (N3810, N2611_t0);
buf BUFF1_888 (N3813, N2607_t0);
buf BUFF1_889 (N3816, N2615_t0);
buf BUFF1_890 (N3819, N2538_t2);
buf BUFF1_891 (N3822, N2546_t2);
buf BUFF1_892 (N3825, N2542_t2);
buf BUFF1_893 (N3828, N2462_t2);
buf BUFF1_894 (N3831, N2550_t2);
buf BUFF1_895 (N3834, N2470_t2);
buf BUFF1_896 (N3837, N2466_t2);
buf BUFF1_897 (N3840, N2478_t2);
buf BUFF1_898 (N3843, N2474_t2);
buf BUFF1_899 (N3846, N2615_t1);
buf BUFF1_900 (N3849, N2611_t1);
buf BUFF1_901 (N3852, N2607_t1);
buf BUFF1_902 (N3855, N2680_t0);
buf BUFF1_903 (N3858, N2729_t2);
buf BUFF1_904 (N3861, N2737_t2);
buf BUFF1_905 (N3864, N2733_t2);
buf BUFF1_906 (N3867, N2745_t2);
buf BUFF1_907 (N3870, N2741_t2);
buf BUFF1_908 (N3873, N2753_t2);
buf BUFF1_909 (N3876, N2749_t2);
buf BUFF1_910 (N3879, N2761_t2);
buf BUFF1_911 (N3882, N2757_t2);
or OR2_912 (N3885, N3033, N2419);
or OR2_913 (N3888, N3032, N2418);
or OR2_914 (N3891, N3020, N2396);
nand NAND2_915 (N3953, N3067_t0, N2117);
not NOT1_916 (N3954, N3067_t1);
nand NAND2_917 (N3955, N3070_t0, N2537);
not NOT1_918 (N3956, N3070_t1);
not NOT1_919 (N3958, N3073_t0);
not NOT1_920 (N3964, N3080_t0);
or OR2_921 (N4193, N1649, N3379);
or OR3_922 (N4303, N1167_t3, N2867, N3130);
not NOT1_923 (N4308, N3061_t0);
not NOT1_924 (N4313, N3064_t0);
nand NAND2_925 (N4326, N2769_t1, N3551);
nand NAND2_926 (N4327, N2766_t1, N3552);
nand NAND2_927 (N4333, N2775_t1, N3569);
nand NAND2_928 (N4334, N2772_t1, N3570);
nand NAND2_929 (N4411, N2787_t1, N3781);
nand NAND2_930 (N4412, N2784_t1, N3782);
nand NAND2_931 (N4463, N3487_t0, N1828);
not NOT1_932 (N4464, N3487_t1);
nand NAND2_933 (N4465, N3490_t0, N1829);
not NOT1_934 (N4466, N3490_t1);
nand NAND2_935 (N4467, N3493_t0, N2267);
not NOT1_936 (N4468, N3493_t1);
nand NAND2_937 (N4469, N3496_t0, N1830);
not NOT1_938 (N4470, N3496_t1);
nand NAND2_939 (N4471, N3499_t0, N1833);
not NOT1_940 (N4472, N3499_t1);
not NOT1_941 (N4473, N3122_t0);
not NOT1_942 (N4474, N3126_t0);
nand NAND2_943 (N4475, N3518_t0, N1840);
not NOT1_944 (N4476, N3518_t1);
nand NAND2_945 (N4477, N3521_t0, N1841);
not NOT1_946 (N4478, N3521_t1);
nand NAND2_947 (N4479, N3524_t0, N2275);
not NOT1_948 (N4480, N3524_t1);
nand NAND2_949 (N4481, N3527_t0, N1842);
not NOT1_950 (N4482, N3527_t1);
nand NAND2_951 (N4483, N3530_t0, N1843);
not NOT1_952 (N4484, N3530_t1);
not NOT1_953 (N4485, N3155_t0);
not NOT1_954 (N4486, N3159_t0);
nand NAND2_955 (N4487, N1721_t1, N3954);
nand NAND2_956 (N4488, N2235_t1, N3956);
not NOT1_957 (N4489, N3535_t0);
nand NAND2_958 (N4490, N3535_t1, N3958);
not NOT1_959 (N4491, N3539_t0);
not NOT1_960 (N4492, N3542_t0);
not NOT1_961 (N4493, N3545_t0);
not NOT1_962 (N4494, N3548_t0);
not NOT1_963 (N4495, N3553_t0);
nand NAND2_964 (N4496, N3553_t1, N3964);
not NOT1_965 (N4497, N3557_t0);
not NOT1_966 (N4498, N3560_t0);
not NOT1_967 (N4499, N3563_t0);
not NOT1_968 (N4500, N3566_t0);
not NOT1_969 (N4501, N3571_t0);
nand NAND2_970 (N4502, N3571_t1, N3167);
not NOT1_971 (N4503, N3574_t0);
not NOT1_972 (N4504, N3577_t0);
not NOT1_973 (N4505, N3580_t0);
not NOT1_974 (N4506, N3583_t0);
nand NAND2_975 (N4507, N3598_t0, N1867);
not NOT1_976 (N4508, N3598_t1);
nand NAND2_977 (N4509, N3601_t0, N1868);
not NOT1_978 (N4510, N3601_t1);
nand NAND2_979 (N4511, N3604_t0, N1869);
not NOT1_980 (N4512, N3604_t1);
nand NAND2_981 (N4513, N3607_t0, N1870);
not NOT1_982 (N4514, N3607_t1);
nand NAND2_983 (N4515, N3610_t0, N1871);
not NOT1_984 (N4516, N3610_t1);
nand NAND2_985 (N4517, N3613_t0, N1872);
not NOT1_986 (N4518, N3613_t1);
nand NAND2_987 (N4519, N3616_t0, N1873);
not NOT1_988 (N4520, N3616_t1);
nand NAND2_989 (N4521, N3619_t0, N1874);
not NOT1_990 (N4522, N3619_t1);
nand NAND2_991 (N4523, N3622_t0, N1875);
not NOT1_992 (N4524, N3622_t1);
nand NAND2_993 (N4525, N3631_t0, N1876);
not NOT1_994 (N4526, N3631_t1);
nand NAND2_995 (N4527, N3634_t0, N1877);
not NOT1_996 (N4528, N3634_t1);
nand NAND2_997 (N4529, N3637_t0, N1878);
not NOT1_998 (N4530, N3637_t1);
nand NAND2_999 (N4531, N3640_t0, N1879);
not NOT1_1000 (N4532, N3640_t1);
nand NAND2_1001 (N4533, N3643_t0, N1880);
not NOT1_1002 (N4534, N3643_t1);
nand NAND2_1003 (N4535, N3646_t0, N1881);
not NOT1_1004 (N4536, N3646_t1);
nand NAND2_1005 (N4537, N3649_t0, N1882);
not NOT1_1006 (N4538, N3649_t1);
nand NAND2_1007 (N4539, N3652_t0, N1883);
not NOT1_1008 (N4540, N3652_t1);
nand NAND2_1009 (N4541, N3655_t0, N1884);
not NOT1_1010 (N4542, N3655_t1);
not NOT1_1011 (N4543, N3658_t0);
and AND2_1012 (N4544, N806_t3, N3293_t0);
and AND2_1013 (N4545, N800_t3, N3287_t0);
and AND2_1014 (N4549, N794_t3, N3281_t0);
and AND2_1015 (N4555, N3273_t0, N786_t3);
and AND2_1016 (N4562, N780_t3, N3267_t0);
and AND2_1017 (N4563, N774_t3, N3355_t0);
and AND2_1018 (N4566, N768_t3, N3349_t0);
and AND2_1019 (N4570, N762_t3, N3343_t0);
not NOT1_1020 (N4575, N3661_t0);
and AND2_1021 (N4576, N806_t4, N3293_t1);
and AND2_1022 (N4577, N800_t4, N3287_t1);
and AND2_1023 (N4581, N794_t4, N3281_t1);
and AND2_1024 (N4586, N786_t4, N3273_t1);
and AND2_1025 (N4592, N780_t4, N3267_t1);
and AND2_1026 (N4593, N774_t4, N3355_t1);
and AND2_1027 (N4597, N768_t4, N3349_t1);
and AND2_1028 (N4603, N762_t4, N3343_t1);
not NOT1_1029 (N4610, N3664_t0);
not NOT1_1030 (N4611, N3667_t0);
not NOT1_1031 (N4612, N3670_t0);
not NOT1_1032 (N4613, N3673_t0);
not NOT1_1033 (N4614, N3676_t0);
not NOT1_1034 (N4615, N3679_t0);
not NOT1_1035 (N4616, N3682_t0);
not NOT1_1036 (N4617, N3685_t0);
not NOT1_1037 (N4618, N3688_t0);
not NOT1_1038 (N4619, N3691_t0);
not NOT1_1039 (N4620, N3694_t0);
not NOT1_1040 (N4621, N3697_t0);
not NOT1_1041 (N4622, N3700_t0);
not NOT1_1042 (N4623, N3703_t0);
not NOT1_1043 (N4624, N3706_t0);
not NOT1_1044 (N4625, N3709_t0);
not NOT1_1045 (N4626, N3712_t0);
not NOT1_1046 (N4627, N3715_t0);
not NOT1_1047 (N4628, N3718_t0);
not NOT1_1048 (N4629, N3721_t0);
and AND2_1049 (N4630, N3448_t0, N2704_t2);
not NOT1_1050 (N4631, N3724_t0);
and AND2_1051 (N4632, N3444_t0, N2700_t2);
not NOT1_1052 (N4633, N3727_t0);
and AND2_1053 (N4634, N3440_t0, N2696_t2);
and AND2_1054 (N4635, N3436_t0, N2692_t2);
not NOT1_1055 (N4636, N3730_t0);
and AND2_1056 (N4637, N3432_t0, N2688_t2);
and AND2_1057 (N4638, N3428_t0, N3311_t0);
and AND2_1058 (N4639, N3424_t0, N3307_t0);
and AND2_1059 (N4640, N3420_t0, N3303_t0);
and AND2_1060 (N4641, N3416_t0, N3299_t0);
not NOT1_1061 (N4642, N3733_t0);
not NOT1_1062 (N4643, N3736_t0);
not NOT1_1063 (N4644, N3739_t0);
not NOT1_1064 (N4645, N3742_t0);
not NOT1_1065 (N4646, N3745_t0);
not NOT1_1066 (N4647, N3748_t0);
not NOT1_1067 (N4648, N3751_t0);
not NOT1_1068 (N4649, N3754_t0);
not NOT1_1069 (N4650, N3757_t0);
not NOT1_1070 (N4651, N3760_t0);
not NOT1_1071 (N4652, N3763_t0);
not NOT1_1072 (N4653, N3375_t0);
and AND2_1073 (N4656, N865_t3, N3410_t0);
and AND2_1074 (N4657, N859_t3, N3404_t0);
and AND2_1075 (N4661, N853_t3, N3398_t0);
and AND2_1076 (N4667, N3390_t0, N845_t3);
and AND2_1077 (N4674, N839_t3, N3384_t0);
and AND2_1078 (N4675, N833_t3, N3334_t0);
and AND2_1079 (N4678, N827_t3, N3328_t0);
and AND2_1080 (N4682, N821_t3, N3322_t0);
and AND2_1081 (N4687, N814_t3, N3315_t0);
not NOT1_1082 (N4693, N3766_t0);
nand NAND2_1083 (N4694, N3766_t1, N3380);
not NOT1_1084 (N4695, N3769_t0);
not NOT1_1085 (N4696, N3772_t0);
not NOT1_1086 (N4697, N3775_t0);
not NOT1_1087 (N4698, N3778_t0);
not NOT1_1088 (N4699, N3783_t0);
not NOT1_1089 (N4700, N3786_t0);
and AND2_1090 (N4701, N865_t4, N3410_t1);
and AND2_1091 (N4702, N859_t4, N3404_t1);
and AND2_1092 (N4706, N853_t4, N3398_t1);
and AND2_1093 (N4711, N845_t4, N3390_t1);
and AND2_1094 (N4717, N839_t4, N3384_t1);
and AND2_1095 (N4718, N833_t4, N3334_t1);
and AND2_1096 (N4722, N827_t4, N3328_t1);
and AND2_1097 (N4728, N821_t4, N3322_t1);
and AND2_1098 (N4735, N814_t4, N3315_t1);
not NOT1_1099 (N4743, N3789_t0);
not NOT1_1100 (N4744, N3792_t0);
not NOT1_1101 (N4745, N3807_t0);
nand NAND2_1102 (N4746, N3807_t1, N3452);
not NOT1_1103 (N4747, N3810_t0);
not NOT1_1104 (N4748, N3813_t0);
not NOT1_1105 (N4749, N3816_t0);
not NOT1_1106 (N4750, N3819_t0);
nand NAND2_1107 (N4751, N3819_t1, N3453);
not NOT1_1108 (N4752, N3822_t0);
not NOT1_1109 (N4753, N3825_t0);
not NOT1_1110 (N4754, N3828_t0);
not NOT1_1111 (N4755, N3831_t0);
and AND2_1112 (N4756, N3482_t0, N3263_t0);
and AND2_1113 (N4757, N3478_t0, N3259_t0);
and AND2_1114 (N4758, N3474_t0, N3255_t0);
and AND2_1115 (N4759, N3470_t0, N3251_t0);
and AND2_1116 (N4760, N3466_t0, N3247_t0);
not NOT1_1117 (N4761, N3846_t0);
and AND2_1118 (N4762, N3462_t0, N2615_t2);
not NOT1_1119 (N4763, N3849_t0);
and AND2_1120 (N4764, N3458_t0, N2611_t2);
not NOT1_1121 (N4765, N3852_t0);
and AND2_1122 (N4766, N3454_t0, N2607_t2);
and AND2_1123 (N4767, N2680_t1, N3381_t0);
not NOT1_1124 (N4768, N3855_t0);
and AND2_1125 (N4769, N3340_t0, N695_t3);
not NOT1_1126 (N4775, N3858_t0);
nand NAND2_1127 (N4776, N3858_t1, N3486);
not NOT1_1128 (N4777, N3861_t0);
not NOT1_1129 (N4778, N3864_t0);
not NOT1_1130 (N4779, N3867_t0);
not NOT1_1131 (N4780, N3870_t0);
not NOT1_1132 (N4781, N3885_t0);
not NOT1_1133 (N4782, N3888_t0);
not NOT1_1134 (N4783, N3891_t0);
or OR2_1135 (N4784, N3131_t0, N3134);
not NOT1_1136 (N4789, N3502_t0);
not NOT1_1137 (N4790, N3131_t1);
not NOT1_1138 (N4793, N3507_t0);
not NOT1_1139 (N4794, N3510_t0);
not NOT1_1140 (N4795, N3515_t0);
buf BUFF1_1141 (N4796, N3114_t0);
not NOT1_1142 (N4799, N3586_t0);
not NOT1_1143 (N4800, N3589_t0);
not NOT1_1144 (N4801, N3592_t0);
not NOT1_1145 (N4802, N3595_t0);
nand NAND2_1146 (N4803, N4326, N4327);
nand NAND2_1147 (N4806, N4333, N4334);
not NOT1_1148 (N4809, N3625_t0);
buf BUFF1_1149 (N4810, N3178_t0);
not NOT1_1150 (N4813, N3628_t0);
buf BUFF1_1151 (N4814, N3202_t0);
buf BUFF1_1152 (N4817, N3221_t0);
buf BUFF1_1153 (N4820, N3293_t2);
buf BUFF1_1154 (N4823, N3287_t2);
buf BUFF1_1155 (N4826, N3281_t2);
buf BUFF1_1156 (N4829, N3273_t2);
buf BUFF1_1157 (N4832, N3267_t2);
buf BUFF1_1158 (N4835, N3355_t2);
buf BUFF1_1159 (N4838, N3349_t2);
buf BUFF1_1160 (N4841, N3343_t2);
nor NOR2_1161 (N4844, N3273_t3, N786_t5);
buf BUFF1_1162 (N4847, N3293_t3);
buf BUFF1_1163 (N4850, N3287_t3);
buf BUFF1_1164 (N4853, N3281_t3);
buf BUFF1_1165 (N4856, N3267_t3);
buf BUFF1_1166 (N4859, N3355_t3);
buf BUFF1_1167 (N4862, N3349_t3);
buf BUFF1_1168 (N4865, N3343_t3);
buf BUFF1_1169 (N4868, N3273_t4);
nor NOR2_1170 (N4871, N786_t6, N3273_t5);
buf BUFF1_1171 (N4874, N3448_t1);
buf BUFF1_1172 (N4877, N3444_t1);
buf BUFF1_1173 (N4880, N3440_t1);
buf BUFF1_1174 (N4883, N3432_t1);
buf BUFF1_1175 (N4886, N3428_t1);
buf BUFF1_1176 (N4889, N3311_t1);
buf BUFF1_1177 (N4892, N3424_t1);
buf BUFF1_1178 (N4895, N3307_t1);
buf BUFF1_1179 (N4898, N3420_t1);
buf BUFF1_1180 (N4901, N3303_t1);
buf BUFF1_1181 (N4904, N3436_t1);
buf BUFF1_1182 (N4907, N3416_t1);
buf BUFF1_1183 (N4910, N3299_t1);
buf BUFF1_1184 (N4913, N3410_t2);
buf BUFF1_1185 (N4916, N3404_t2);
buf BUFF1_1186 (N4919, N3398_t2);
buf BUFF1_1187 (N4922, N3390_t2);
buf BUFF1_1188 (N4925, N3384_t2);
buf BUFF1_1189 (N4928, N3334_t2);
buf BUFF1_1190 (N4931, N3328_t2);
buf BUFF1_1191 (N4934, N3322_t2);
buf BUFF1_1192 (N4937, N3315_t2);
nor NOR2_1193 (N4940, N3390_t3, N845_t5);
buf BUFF1_1194 (N4943, N3315_t3);
buf BUFF1_1195 (N4946, N3328_t3);
buf BUFF1_1196 (N4949, N3322_t3);
buf BUFF1_1197 (N4952, N3384_t3);
buf BUFF1_1198 (N4955, N3334_t3);
buf BUFF1_1199 (N4958, N3398_t3);
buf BUFF1_1200 (N4961, N3390_t4);
buf BUFF1_1201 (N4964, N3410_t3);
buf BUFF1_1202 (N4967, N3404_t3);
buf BUFF1_1203 (N4970, N3340_t1);
buf BUFF1_1204 (N4973, N3349_t4);
buf BUFF1_1205 (N4976, N3343_t4);
buf BUFF1_1206 (N4979, N3267_t4);
buf BUFF1_1207 (N4982, N3355_t4);
buf BUFF1_1208 (N4985, N3281_t4);
buf BUFF1_1209 (N4988, N3273_t6);
buf BUFF1_1210 (N4991, N3293_t4);
buf BUFF1_1211 (N4994, N3287_t4);
nand NAND2_1212 (N4997, N4411, N4412);
buf BUFF1_1213 (N5000, N3410_t4);
buf BUFF1_1214 (N5003, N3404_t4);
buf BUFF1_1215 (N5006, N3398_t4);
buf BUFF1_1216 (N5009, N3384_t4);
buf BUFF1_1217 (N5012, N3334_t4);
buf BUFF1_1218 (N5015, N3328_t4);
buf BUFF1_1219 (N5018, N3322_t4);
buf BUFF1_1220 (N5021, N3390_t5);
buf BUFF1_1221 (N5024, N3315_t4);
nor NOR2_1222 (N5027, N845_t6, N3390_t6);
nor NOR2_1223 (N5030, N814_t5, N3315_t5);
buf BUFF1_1224 (N5033, N3299_t2);
buf BUFF1_1225 (N5036, N3307_t2);
buf BUFF1_1226 (N5039, N3303_t2);
buf BUFF1_1227 (N5042, N3311_t2);
not NOT1_1228 (N5045, N3795_t0);
not NOT1_1229 (N5046, N3798_t0);
not NOT1_1230 (N5047, N3801_t0);
not NOT1_1231 (N5048, N3804_t0);
buf BUFF1_1232 (N5049, N3247_t1);
buf BUFF1_1233 (N5052, N3255_t1);
buf BUFF1_1234 (N5055, N3251_t1);
buf BUFF1_1235 (N5058, N3263_t1);
buf BUFF1_1236 (N5061, N3259_t1);
not NOT1_1237 (N5064, N3834_t0);
not NOT1_1238 (N5065, N3837_t0);
not NOT1_1239 (N5066, N3840_t0);
not NOT1_1240 (N5067, N3843_t0);
buf BUFF1_1241 (N5068, N3482_t1);
buf BUFF1_1242 (N5071, N3263_t2);
buf BUFF1_1243 (N5074, N3478_t1);
buf BUFF1_1244 (N5077, N3259_t2);
buf BUFF1_1245 (N5080, N3474_t1);
buf BUFF1_1246 (N5083, N3255_t2);
buf BUFF1_1247 (N5086, N3466_t1);
buf BUFF1_1248 (N5089, N3247_t2);
buf BUFF1_1249 (N5092, N3462_t1);
buf BUFF1_1250 (N5095, N3458_t1);
buf BUFF1_1251 (N5098, N3454_t1);
buf BUFF1_1252 (N5101, N3470_t1);
buf BUFF1_1253 (N5104, N3251_t2);
buf BUFF1_1254 (N5107, N3381_t1);
not NOT1_1255 (N5110, N3873_t0);
not NOT1_1256 (N5111, N3876_t0);
not NOT1_1257 (N5112, N3879_t0);
not NOT1_1258 (N5113, N3882_t0);
buf BUFF1_1259 (N5114, N3458_t2);
buf BUFF1_1260 (N5117, N3454_t2);
buf BUFF1_1261 (N5120, N3466_t2);
buf BUFF1_1262 (N5123, N3462_t2);
buf BUFF1_1263 (N5126, N3474_t2);
buf BUFF1_1264 (N5129, N3470_t2);
buf BUFF1_1265 (N5132, N3482_t2);
buf BUFF1_1266 (N5135, N3478_t2);
buf BUFF1_1267 (N5138, N3416_t2);
buf BUFF1_1268 (N5141, N3424_t2);
buf BUFF1_1269 (N5144, N3420_t2);
buf BUFF1_1270 (N5147, N3432_t2);
buf BUFF1_1271 (N5150, N3428_t2);
buf BUFF1_1272 (N5153, N3440_t2);
buf BUFF1_1273 (N5156, N3436_t2);
buf BUFF1_1274 (N5159, N3448_t2);
buf BUFF1_1275 (N5162, N3444_t2);
nand NAND2_1276 (N5165, N4486, N4485);
nand NAND2_1277 (N5166, N4474, N4473);
nand NAND2_1278 (N5167, N1290_t1, N4464);
nand NAND2_1279 (N5168, N1293_t1, N4466);
nand NAND2_1280 (N5169, N2074_t1, N4468);
nand NAND2_1281 (N5170, N1296_t1, N4470);
nand NAND2_1282 (N5171, N1302_t1, N4472);
nand NAND2_1283 (N5172, N1314_t1, N4476);
nand NAND2_1284 (N5173, N1317_t1, N4478);
nand NAND2_1285 (N5174, N2081_t1, N4480);
nand NAND2_1286 (N5175, N1320_t1, N4482);
nand NAND2_1287 (N5176, N1323_t1, N4484);
nand NAND2_1288 (N5177, N3953, N4487);
nand NAND2_1289 (N5178, N3955, N4488);
nand NAND2_1290 (N5179, N3073_t1, N4489);
nand NAND2_1291 (N5180, N3542_t1, N4491);
nand NAND2_1292 (N5181, N3539_t1, N4492);
nand NAND2_1293 (N5182, N3548_t1, N4493);
nand NAND2_1294 (N5183, N3545_t1, N4494);
nand NAND2_1295 (N5184, N3080_t1, N4495);
nand NAND2_1296 (N5185, N3560_t1, N4497);
nand NAND2_1297 (N5186, N3557_t1, N4498);
nand NAND2_1298 (N5187, N3566_t1, N4499);
nand NAND2_1299 (N5188, N3563_t1, N4500);
nand NAND2_1300 (N5189, N2778_t1, N4501);
nand NAND2_1301 (N5190, N3577_t1, N4503);
nand NAND2_1302 (N5191, N3574_t1, N4504);
nand NAND2_1303 (N5192, N3583_t1, N4505);
nand NAND2_1304 (N5193, N3580_t1, N4506);
nand NAND2_1305 (N5196, N1326_t1, N4508);
nand NAND2_1306 (N5197, N1329_t1, N4510);
nand NAND2_1307 (N5198, N1332_t1, N4512);
nand NAND2_1308 (N5199, N1335_t1, N4514);
nand NAND2_1309 (N5200, N1338_t1, N4516);
nand NAND2_1310 (N5201, N1341_t1, N4518);
nand NAND2_1311 (N5202, N1344_t1, N4520);
nand NAND2_1312 (N5203, N1347_t1, N4522);
nand NAND2_1313 (N5204, N1350_t1, N4524);
nand NAND2_1314 (N5205, N1353_t1, N4526);
nand NAND2_1315 (N5206, N1356_t1, N4528);
nand NAND2_1316 (N5207, N1359_t1, N4530);
nand NAND2_1317 (N5208, N1362_t1, N4532);
nand NAND2_1318 (N5209, N1365_t1, N4534);
nand NAND2_1319 (N5210, N1368_t1, N4536);
nand NAND2_1320 (N5211, N1371_t1, N4538);
nand NAND2_1321 (N5212, N1374_t1, N4540);
nand NAND2_1322 (N5213, N1377_t1, N4542);
nand NAND2_1323 (N5283, N3670_t1, N4611);
nand NAND2_1324 (N5284, N3667_t1, N4612);
nand NAND2_1325 (N5285, N3676_t1, N4613);
nand NAND2_1326 (N5286, N3673_t1, N4614);
nand NAND2_1327 (N5287, N3682_t1, N4615);
nand NAND2_1328 (N5288, N3679_t1, N4616);
nand NAND2_1329 (N5289, N3688_t1, N4617);
nand NAND2_1330 (N5290, N3685_t1, N4618);
nand NAND2_1331 (N5291, N3694_t1, N4619);
nand NAND2_1332 (N5292, N3691_t1, N4620);
nand NAND2_1333 (N5293, N3700_t1, N4621);
nand NAND2_1334 (N5294, N3697_t1, N4622);
nand NAND2_1335 (N5295, N3706_t1, N4623);
nand NAND2_1336 (N5296, N3703_t1, N4624);
nand NAND2_1337 (N5297, N3712_t1, N4625);
nand NAND2_1338 (N5298, N3709_t1, N4626);
nand NAND2_1339 (N5299, N3718_t1, N4627);
nand NAND2_1340 (N5300, N3715_t1, N4628);
nand NAND2_1341 (N5314, N3739_t1, N4643);
nand NAND2_1342 (N5315, N3736_t1, N4644);
nand NAND2_1343 (N5316, N3745_t1, N4645);
nand NAND2_1344 (N5317, N3742_t1, N4646);
nand NAND2_1345 (N5318, N3751_t1, N4647);
nand NAND2_1346 (N5319, N3748_t1, N4648);
nand NAND2_1347 (N5320, N3757_t1, N4649);
nand NAND2_1348 (N5321, N3754_t1, N4650);
nand NAND2_1349 (N5322, N3763_t1, N4651);
nand NAND2_1350 (N5323, N3760_t1, N4652);
not NOT1_1351 (N5324, N4193_t0);
nand NAND2_1352 (N5363, N2781_t1, N4693);
nand NAND2_1353 (N5364, N3772_t1, N4695);
nand NAND2_1354 (N5365, N3769_t1, N4696);
nand NAND2_1355 (N5366, N3778_t1, N4697);
nand NAND2_1356 (N5367, N3775_t1, N4698);
nand NAND2_1357 (N5425, N2790_t1, N4745);
nand NAND2_1358 (N5426, N3813_t1, N4747);
nand NAND2_1359 (N5427, N3810_t1, N4748);
nand NAND2_1360 (N5429, N2793_t1, N4750);
nand NAND2_1361 (N5430, N3825_t1, N4752);
nand NAND2_1362 (N5431, N3822_t1, N4753);
nand NAND2_1363 (N5432, N3831_t1, N4754);
nand NAND2_1364 (N5433, N3828_t1, N4755);
nand NAND2_1365 (N5451, N2796_t1, N4775);
nand NAND2_1366 (N5452, N3864_t1, N4777);
nand NAND2_1367 (N5453, N3861_t1, N4778);
nand NAND2_1368 (N5454, N3870_t1, N4779);
nand NAND2_1369 (N5455, N3867_t1, N4780);
nand NAND2_1370 (N5456, N3888_t1, N4781);
nand NAND2_1371 (N5457, N3885_t1, N4782);
not NOT1_1372 (N5469, N4303_t0);
nand NAND2_1373 (N5474, N3589_t1, N4799);
nand NAND2_1374 (N5475, N3586_t1, N4800);
nand NAND2_1375 (N5476, N3595_t1, N4801);
nand NAND2_1376 (N5477, N3592_t1, N4802);
nand NAND2_1377 (N5571, N3798_t1, N5045);
nand NAND2_1378 (N5572, N3795_t1, N5046);
nand NAND2_1379 (N5573, N3804_t1, N5047);
nand NAND2_1380 (N5574, N3801_t1, N5048);
nand NAND2_1381 (N5584, N3837_t1, N5064);
nand NAND2_1382 (N5585, N3834_t1, N5065);
nand NAND2_1383 (N5586, N3843_t1, N5066);
nand NAND2_1384 (N5587, N3840_t1, N5067);
nand NAND2_1385 (N5602, N3876_t1, N5110);
nand NAND2_1386 (N5603, N3873_t1, N5111);
nand NAND2_1387 (N5604, N3882_t1, N5112);
nand NAND2_1388 (N5605, N3879_t1, N5113);
nand NAND2_1389 (N5631, N5324, N4653);
nand NAND2_1390 (N5632, N4463, N5167);
nand NAND2_1391 (N5640, N4465, N5168);
nand NAND2_1392 (N5654, N4467, N5169);
nand NAND2_1393 (N5670, N4469, N5170);
nand NAND2_1394 (N5683, N4471, N5171);
nand NAND2_1395 (N5690, N4475, N5172);
nand NAND2_1396 (N5697, N4477, N5173);
nand NAND2_1397 (N5707, N4479, N5174);
nand NAND2_1398 (N5718, N4481, N5175);
nand NAND2_1399 (N5728, N4483, N5176);
not NOT1_1400 (N5735, N5177);
nand NAND2_1401 (N5736, N5179, N4490);
nand NAND2_1402 (N5740, N5180, N5181);
nand NAND2_1403 (N5744, N5182, N5183);
nand NAND2_1404 (N5747, N5184, N4496);
nand NAND2_1405 (N5751, N5185, N5186);
nand NAND2_1406 (N5755, N5187, N5188);
nand NAND2_1407 (N5758, N5189, N4502);
nand NAND2_1408 (N5762, N5190, N5191);
nand NAND2_1409 (N5766, N5192, N5193);
not NOT1_1410 (N5769, N4803_t0);
not NOT1_1411 (N5770, N4806_t0);
nand NAND2_1412 (N5771, N4507, N5196);
nand NAND2_1413 (N5778, N4509, N5197);
nand NAND2_1414 (N5789, N4511, N5198);
nand NAND2_1415 (N5799, N4513, N5199);
nand NAND2_1416 (N5807, N4515, N5200);
nand NAND2_1417 (N5821, N4517, N5201);
nand NAND2_1418 (N5837, N4519, N5202);
nand NAND2_1419 (N5850, N4521, N5203);
nand NAND2_1420 (N5856, N4523, N5204);
nand NAND2_1421 (N5863, N4525, N5205);
nand NAND2_1422 (N5870, N4527, N5206);
nand NAND2_1423 (N5881, N4529, N5207);
nand NAND2_1424 (N5892, N4531, N5208);
nand NAND2_1425 (N5898, N4533, N5209);
nand NAND2_1426 (N5905, N4535, N5210);
nand NAND2_1427 (N5915, N4537, N5211);
nand NAND2_1428 (N5926, N4539, N5212);
nand NAND2_1429 (N5936, N4541, N5213);
not NOT1_1430 (N5943, N4817_t0);
nand NAND2_1431 (N5944, N4820_t0, N1931);
not NOT1_1432 (N5945, N4820_t1);
nand NAND2_1433 (N5946, N4823_t0, N1932);
not NOT1_1434 (N5947, N4823_t1);
nand NAND2_1435 (N5948, N4826_t0, N1933);
not NOT1_1436 (N5949, N4826_t1);
nand NAND2_1437 (N5950, N4829_t0, N1934);
not NOT1_1438 (N5951, N4829_t1);
nand NAND2_1439 (N5952, N4832_t0, N1935);
not NOT1_1440 (N5953, N4832_t1);
nand NAND2_1441 (N5954, N4835_t0, N1936);
not NOT1_1442 (N5955, N4835_t1);
nand NAND2_1443 (N5956, N4838_t0, N1937);
not NOT1_1444 (N5957, N4838_t1);
nand NAND2_1445 (N5958, N4841_t0, N1938);
not NOT1_1446 (N5959, N4841_t1);
and AND2_1447 (N5960, N2674_t2, N4769_t0);
not NOT1_1448 (N5966, N4844_t0);
nand NAND2_1449 (N5967, N4847_t0, N1939);
not NOT1_1450 (N5968, N4847_t1);
nand NAND2_1451 (N5969, N4850_t0, N1940);
not NOT1_1452 (N5970, N4850_t1);
nand NAND2_1453 (N5971, N4853_t0, N1941);
not NOT1_1454 (N5972, N4853_t1);
nand NAND2_1455 (N5973, N4856_t0, N1942);
not NOT1_1456 (N5974, N4856_t1);
nand NAND2_1457 (N5975, N4859_t0, N1943);
not NOT1_1458 (N5976, N4859_t1);
nand NAND2_1459 (N5977, N4862_t0, N1944);
not NOT1_1460 (N5978, N4862_t1);
nand NAND2_1461 (N5979, N4865_t0, N1945);
not NOT1_1462 (N5980, N4865_t1);
and AND2_1463 (N5981, N2674_t3, N4769_t1);
nand NAND2_1464 (N5989, N4868_t0, N1946);
not NOT1_1465 (N5990, N4868_t1);
nand NAND2_1466 (N5991, N5283, N5284);
nand NAND2_1467 (N5996, N5285, N5286);
nand NAND2_1468 (N6000, N5287, N5288);
nand NAND2_1469 (N6003, N5289, N5290);
nand NAND2_1470 (N6009, N5291, N5292);
nand NAND2_1471 (N6014, N5293, N5294);
nand NAND2_1472 (N6018, N5295, N5296);
nand NAND2_1473 (N6021, N5297, N5298);
nand NAND2_1474 (N6022, N5299, N5300);
not NOT1_1475 (N6023, N4874_t0);
nand NAND2_1476 (N6024, N4874_t1, N4629);
not NOT1_1477 (N6025, N4877_t0);
nand NAND2_1478 (N6026, N4877_t1, N4631);
not NOT1_1479 (N6027, N4880_t0);
nand NAND2_1480 (N6028, N4880_t1, N4633);
not NOT1_1481 (N6029, N4883_t0);
nand NAND2_1482 (N6030, N4883_t1, N4636);
not NOT1_1483 (N6031, N4886_t0);
not NOT1_1484 (N6032, N4889_t0);
not NOT1_1485 (N6033, N4892_t0);
not NOT1_1486 (N6034, N4895_t0);
not NOT1_1487 (N6035, N4898_t0);
not NOT1_1488 (N6036, N4901_t0);
not NOT1_1489 (N6037, N4904_t0);
nand NAND2_1490 (N6038, N4904_t1, N4642);
not NOT1_1491 (N6039, N4907_t0);
not NOT1_1492 (N6040, N4910_t0);
nand NAND2_1493 (N6041, N5314, N5315);
nand NAND2_1494 (N6047, N5316, N5317);
nand NAND2_1495 (N6052, N5318, N5319);
nand NAND2_1496 (N6056, N5320, N5321);
nand NAND2_1497 (N6059, N5322, N5323);
nand NAND2_1498 (N6060, N4913_t0, N1968);
not NOT1_1499 (N6061, N4913_t1);
nand NAND2_1500 (N6062, N4916_t0, N1969);
not NOT1_1501 (N6063, N4916_t1);
nand NAND2_1502 (N6064, N4919_t0, N1970);
not NOT1_1503 (N6065, N4919_t1);
nand NAND2_1504 (N6066, N4922_t0, N1971);
not NOT1_1505 (N6067, N4922_t1);
nand NAND2_1506 (N6068, N4925_t0, N1972);
not NOT1_1507 (N6069, N4925_t1);
nand NAND2_1508 (N6070, N4928_t0, N1973);
not NOT1_1509 (N6071, N4928_t1);
nand NAND2_1510 (N6072, N4931_t0, N1974);
not NOT1_1511 (N6073, N4931_t1);
nand NAND2_1512 (N6074, N4934_t0, N1975);
not NOT1_1513 (N6075, N4934_t1);
nand NAND2_1514 (N6076, N4937_t0, N1976);
not NOT1_1515 (N6077, N4937_t1);
not NOT1_1516 (N6078, N4940_t0);
nand NAND2_1517 (N6079, N5363, N4694);
nand NAND2_1518 (N6083, N5364, N5365);
nand NAND2_1519 (N6087, N5366, N5367);
not NOT1_1520 (N6090, N4943_t0);
nand NAND2_1521 (N6091, N4943_t1, N4699);
not NOT1_1522 (N6092, N4946_t0);
not NOT1_1523 (N6093, N4949_t0);
not NOT1_1524 (N6094, N4952_t0);
not NOT1_1525 (N6095, N4955_t0);
not NOT1_1526 (N6096, N4970_t0);
nand NAND2_1527 (N6097, N4970_t1, N4700);
not NOT1_1528 (N6098, N4973_t0);
not NOT1_1529 (N6099, N4976_t0);
not NOT1_1530 (N6100, N4979_t0);
not NOT1_1531 (N6101, N4982_t0);
not NOT1_1532 (N6102, N4997_t0);
nand NAND2_1533 (N6103, N5000_t0, N2015);
not NOT1_1534 (N6104, N5000_t1);
nand NAND2_1535 (N6105, N5003_t0, N2016);
not NOT1_1536 (N6106, N5003_t1);
nand NAND2_1537 (N6107, N5006_t0, N2017);
not NOT1_1538 (N6108, N5006_t1);
nand NAND2_1539 (N6109, N5009_t0, N2018);
not NOT1_1540 (N6110, N5009_t1);
nand NAND2_1541 (N6111, N5012_t0, N2019);
not NOT1_1542 (N6112, N5012_t1);
nand NAND2_1543 (N6113, N5015_t0, N2020);
not NOT1_1544 (N6114, N5015_t1);
nand NAND2_1545 (N6115, N5018_t0, N2021);
not NOT1_1546 (N6116, N5018_t1);
nand NAND2_1547 (N6117, N5021_t0, N2022);
not NOT1_1548 (N6118, N5021_t1);
nand NAND2_1549 (N6119, N5024_t0, N2023);
not NOT1_1550 (N6120, N5024_t1);
not NOT1_1551 (N6121, N5033_t0);
nand NAND2_1552 (N6122, N5033_t1, N4743);
not NOT1_1553 (N6123, N5036_t0);
not NOT1_1554 (N6124, N5039_t0);
nand NAND2_1555 (N6125, N5042_t0, N4744);
not NOT1_1556 (N6126, N5042_t1);
nand NAND2_1557 (N6127, N5425, N4746);
nand NAND2_1558 (N6131, N5426, N5427);
not NOT1_1559 (N6135, N5049_t0);
nand NAND2_1560 (N6136, N5049_t1, N4749);
nand NAND2_1561 (N6137, N5429, N4751);
nand NAND2_1562 (N6141, N5430, N5431);
nand NAND2_1563 (N6145, N5432, N5433);
not NOT1_1564 (N6148, N5068_t0);
not NOT1_1565 (N6149, N5071_t0);
not NOT1_1566 (N6150, N5074_t0);
not NOT1_1567 (N6151, N5077_t0);
not NOT1_1568 (N6152, N5080_t0);
not NOT1_1569 (N6153, N5083_t0);
not NOT1_1570 (N6154, N5086_t0);
not NOT1_1571 (N6155, N5089_t0);
not NOT1_1572 (N6156, N5092_t0);
nand NAND2_1573 (N6157, N5092_t1, N4761);
not NOT1_1574 (N6158, N5095_t0);
nand NAND2_1575 (N6159, N5095_t1, N4763);
not NOT1_1576 (N6160, N5098_t0);
nand NAND2_1577 (N6161, N5098_t1, N4765);
not NOT1_1578 (N6162, N5101_t0);
not NOT1_1579 (N6163, N5104_t0);
nand NAND2_1580 (N6164, N5107_t0, N4768);
not NOT1_1581 (N6165, N5107_t1);
nand NAND2_1582 (N6166, N5451, N4776);
nand NAND2_1583 (N6170, N5452, N5453);
nand NAND2_1584 (N6174, N5454, N5455);
nand NAND2_1585 (N6177, N5456, N5457);
not NOT1_1586 (N6181, N5114_t0);
not NOT1_1587 (N6182, N5117_t0);
not NOT1_1588 (N6183, N5120_t0);
not NOT1_1589 (N6184, N5123_t0);
not NOT1_1590 (N6185, N5138_t0);
nand NAND2_1591 (N6186, N5138_t1, N4783);
not NOT1_1592 (N6187, N5141_t0);
not NOT1_1593 (N6188, N5144_t0);
not NOT1_1594 (N6189, N5147_t0);
not NOT1_1595 (N6190, N5150_t0);
not NOT1_1596 (N6191, N4784_t0);
nand NAND2_1597 (N6192, N4784_t1, N2230);
not NOT1_1598 (N6193, N4790_t0);
nand NAND2_1599 (N6194, N4790_t1, N2765);
not NOT1_1600 (N6195, N4796_t0);
nand NAND2_1601 (N6196, N5476, N5477);
nand NAND2_1602 (N6199, N5474, N5475);
not NOT1_1603 (N6202, N4810_t0);
not NOT1_1604 (N6203, N4814_t0);
buf BUFF1_1605 (N6204, N4769_t2);
buf BUFF1_1606 (N6207, N4555_t0);
buf BUFF1_1607 (N6210, N4769_t3);
not NOT1_1608 (N6213, N4871_t0);
buf BUFF1_1609 (N6214, N4586_t0);
nor NOR2_1610 (N6217, N2674_t4, N4769_t4);
buf BUFF1_1611 (N6220, N4667_t0);
not NOT1_1612 (N6223, N4958_t0);
not NOT1_1613 (N6224, N4961_t0);
not NOT1_1614 (N6225, N4964_t0);
not NOT1_1615 (N6226, N4967_t0);
not NOT1_1616 (N6227, N4985_t0);
not NOT1_1617 (N6228, N4988_t0);
not NOT1_1618 (N6229, N4991_t0);
not NOT1_1619 (N6230, N4994_t0);
not NOT1_1620 (N6231, N5027_t0);
buf BUFF1_1621 (N6232, N4711_t0);
not NOT1_1622 (N6235, N5030_t0);
buf BUFF1_1623 (N6236, N4735_t0);
not NOT1_1624 (N6239, N5052_t0);
not NOT1_1625 (N6240, N5055_t0);
not NOT1_1626 (N6241, N5058_t0);
not NOT1_1627 (N6242, N5061_t0);
nand NAND2_1628 (N6243, N5573, N5574);
nand NAND2_1629 (N6246, N5571, N5572);
nand NAND2_1630 (N6249, N5586, N5587);
nand NAND2_1631 (N6252, N5584, N5585);
not NOT1_1632 (N6255, N5126_t0);
not NOT1_1633 (N6256, N5129_t0);
not NOT1_1634 (N6257, N5132_t0);
not NOT1_1635 (N6258, N5135_t0);
not NOT1_1636 (N6259, N5153_t0);
not NOT1_1637 (N6260, N5156_t0);
not NOT1_1638 (N6261, N5159_t0);
not NOT1_1639 (N6262, N5162_t0);
nand NAND2_1640 (N6263, N5604, N5605);
nand NAND2_1641 (N6266, N5602, N5603);
nand NAND2_1642 (N6540, N1380_t1, N5945);
nand NAND2_1643 (N6541, N1383_t1, N5947);
nand NAND2_1644 (N6542, N1386_t1, N5949);
nand NAND2_1645 (N6543, N1389_t1, N5951);
nand NAND2_1646 (N6544, N1392_t1, N5953);
nand NAND2_1647 (N6545, N1395_t1, N5955);
nand NAND2_1648 (N6546, N1398_t1, N5957);
nand NAND2_1649 (N6547, N1401_t1, N5959);
nand NAND2_1650 (N6555, N1404_t1, N5968);
nand NAND2_1651 (N6556, N1407_t1, N5970);
nand NAND2_1652 (N6557, N1410_t1, N5972);
nand NAND2_1653 (N6558, N1413_t1, N5974);
nand NAND2_1654 (N6559, N1416_t1, N5976);
nand NAND2_1655 (N6560, N1419_t1, N5978);
nand NAND2_1656 (N6561, N1422_t1, N5980);
nand NAND2_1657 (N6569, N1425_t1, N5990);
nand NAND2_1658 (N6594, N3721_t1, N6023);
nand NAND2_1659 (N6595, N3724_t1, N6025);
nand NAND2_1660 (N6596, N3727_t1, N6027);
nand NAND2_1661 (N6597, N3730_t1, N6029);
nand NAND2_1662 (N6598, N4889_t1, N6031);
nand NAND2_1663 (N6599, N4886_t1, N6032);
nand NAND2_1664 (N6600, N4895_t1, N6033);
nand NAND2_1665 (N6601, N4892_t1, N6034);
nand NAND2_1666 (N6602, N4901_t1, N6035);
nand NAND2_1667 (N6603, N4898_t1, N6036);
nand NAND2_1668 (N6604, N3733_t1, N6037);
nand NAND2_1669 (N6605, N4910_t1, N6039);
nand NAND2_1670 (N6606, N4907_t1, N6040);
nand NAND2_1671 (N6621, N1434_t1, N6061);
nand NAND2_1672 (N6622, N1437_t1, N6063);
nand NAND2_1673 (N6623, N1440_t1, N6065);
nand NAND2_1674 (N6624, N1443_t1, N6067);
nand NAND2_1675 (N6625, N1446_t1, N6069);
nand NAND2_1676 (N6626, N1449_t1, N6071);
nand NAND2_1677 (N6627, N1452_t1, N6073);
nand NAND2_1678 (N6628, N1455_t1, N6075);
nand NAND2_1679 (N6629, N1458_t1, N6077);
nand NAND2_1680 (N6639, N3783_t1, N6090);
nand NAND2_1681 (N6640, N4949_t1, N6092);
nand NAND2_1682 (N6641, N4946_t1, N6093);
nand NAND2_1683 (N6642, N4955_t1, N6094);
nand NAND2_1684 (N6643, N4952_t1, N6095);
nand NAND2_1685 (N6644, N3786_t1, N6096);
nand NAND2_1686 (N6645, N4976_t1, N6098);
nand NAND2_1687 (N6646, N4973_t1, N6099);
nand NAND2_1688 (N6647, N4982_t1, N6100);
nand NAND2_1689 (N6648, N4979_t1, N6101);
nand NAND2_1690 (N6649, N1461_t1, N6104);
nand NAND2_1691 (N6650, N1464_t1, N6106);
nand NAND2_1692 (N6651, N1467_t1, N6108);
nand NAND2_1693 (N6652, N1470_t1, N6110);
nand NAND2_1694 (N6653, N1473_t1, N6112);
nand NAND2_1695 (N6654, N1476_t1, N6114);
nand NAND2_1696 (N6655, N1479_t1, N6116);
nand NAND2_1697 (N6656, N1482_t1, N6118);
nand NAND2_1698 (N6657, N1485_t1, N6120);
nand NAND2_1699 (N6658, N3789_t1, N6121);
nand NAND2_1700 (N6659, N5039_t1, N6123);
nand NAND2_1701 (N6660, N5036_t1, N6124);
nand NAND2_1702 (N6661, N3792_t1, N6126);
nand NAND2_1703 (N6668, N3816_t1, N6135);
nand NAND2_1704 (N6677, N5071_t1, N6148);
nand NAND2_1705 (N6678, N5068_t1, N6149);
nand NAND2_1706 (N6679, N5077_t1, N6150);
nand NAND2_1707 (N6680, N5074_t1, N6151);
nand NAND2_1708 (N6681, N5083_t1, N6152);
nand NAND2_1709 (N6682, N5080_t1, N6153);
nand NAND2_1710 (N6683, N5089_t1, N6154);
nand NAND2_1711 (N6684, N5086_t1, N6155);
nand NAND2_1712 (N6685, N3846_t1, N6156);
nand NAND2_1713 (N6686, N3849_t1, N6158);
nand NAND2_1714 (N6687, N3852_t1, N6160);
nand NAND2_1715 (N6688, N5104_t1, N6162);
nand NAND2_1716 (N6689, N5101_t1, N6163);
nand NAND2_1717 (N6690, N3855_t1, N6165);
nand NAND2_1718 (N6702, N5117_t1, N6181);
nand NAND2_1719 (N6703, N5114_t1, N6182);
nand NAND2_1720 (N6704, N5123_t1, N6183);
nand NAND2_1721 (N6705, N5120_t1, N6184);
nand NAND2_1722 (N6706, N3891_t1, N6185);
nand NAND2_1723 (N6707, N5144_t1, N6187);
nand NAND2_1724 (N6708, N5141_t1, N6188);
nand NAND2_1725 (N6709, N5150_t1, N6189);
nand NAND2_1726 (N6710, N5147_t1, N6190);
nand NAND2_1727 (N6711, N1708_t1, N6191);
nand NAND2_1728 (N6712, N2231_t1, N6193);
nand NAND2_1729 (N6729, N4961_t1, N6223);
nand NAND2_1730 (N6730, N4958_t1, N6224);
nand NAND2_1731 (N6731, N4967_t1, N6225);
nand NAND2_1732 (N6732, N4964_t1, N6226);
nand NAND2_1733 (N6733, N4988_t1, N6227);
nand NAND2_1734 (N6734, N4985_t1, N6228);
nand NAND2_1735 (N6735, N4994_t1, N6229);
nand NAND2_1736 (N6736, N4991_t1, N6230);
nand NAND2_1737 (N6741, N5055_t1, N6239);
nand NAND2_1738 (N6742, N5052_t1, N6240);
nand NAND2_1739 (N6743, N5061_t1, N6241);
nand NAND2_1740 (N6744, N5058_t1, N6242);
nand NAND2_1741 (N6751, N5129_t1, N6255);
nand NAND2_1742 (N6752, N5126_t1, N6256);
nand NAND2_1743 (N6753, N5135_t1, N6257);
nand NAND2_1744 (N6754, N5132_t1, N6258);
nand NAND2_1745 (N6755, N5156_t1, N6259);
nand NAND2_1746 (N6756, N5153_t1, N6260);
nand NAND2_1747 (N6757, N5162_t1, N6261);
nand NAND2_1748 (N6758, N5159_t1, N6262);
not NOT1_1749 (N6761, N5892_t0);
and AND5_1750 (N6762, N5683_t0, N5670_t0, N5654_t0, N5640_t0, N5632_t0);
and AND2_1751 (N6766, N5632_t1, N3097_t0);
and AND3_1752 (N6767, N5640_t1, N5632_t2, N3101_t0);
and AND4_1753 (N6768, N5654_t1, N5632_t3, N3107_t0, N5640_t2);
and AND5_1754 (N6769, N5670_t1, N5654_t2, N5632_t4, N3114_t1, N5640_t3);
and AND2_1755 (N6770, N5640_t4, N3101_t1);
and AND3_1756 (N6771, N5654_t3, N3107_t1, N5640_t5);
and AND4_1757 (N6772, N5670_t2, N5654_t4, N3114_t2, N5640_t6);
and AND4_1758 (N6773, N5683_t1, N5654_t5, N5640_t7, N5670_t3);
and AND2_1759 (N6774, N5640_t8, N3101_t2);
and AND3_1760 (N6775, N5654_t6, N3107_t2, N5640_t9);
and AND4_1761 (N6776, N5670_t4, N5654_t7, N3114_t3, N5640_t10);
and AND2_1762 (N6777, N5654_t8, N3107_t3);
and AND3_1763 (N6778, N5670_t5, N5654_t9, N3114_t4);
and AND3_1764 (N6779, N5683_t2, N5654_t10, N5670_t6);
and AND2_1765 (N6780, N5654_t11, N3107_t4);
and AND3_1766 (N6781, N5670_t7, N5654_t12, N3114_t5);
and AND2_1767 (N6782, N5670_t8, N3114_t6);
and AND2_1768 (N6783, N5683_t3, N5670_t9);
and AND5_1769 (N6784, N5697_t0, N5728_t0, N5707_t0, N5690_t0, N5718_t0);
and AND2_1770 (N6787, N5690_t1, N3137_t0);
and AND3_1771 (N6788, N5697_t1, N5690_t2, N3140_t0);
and AND4_1772 (N6789, N5707_t1, N5690_t3, N3144_t0, N5697_t2);
and AND5_1773 (N6790, N5718_t1, N5707_t2, N5690_t4, N3149_t0, N5697_t3);
and AND2_1774 (N6791, N5697_t4, N3140_t1);
and AND3_1775 (N6792, N5707_t3, N3144_t1, N5697_t5);
and AND4_1776 (N6793, N5718_t2, N5707_t4, N3149_t1, N5697_t6);
and AND2_1777 (N6794, N3144_t2, N5707_t5);
and AND3_1778 (N6795, N5718_t3, N5707_t6, N3149_t2);
and AND2_1779 (N6796, N5718_t4, N3149_t3);
not NOT1_1780 (N6797, N5736_t0);
not NOT1_1781 (N6800, N5740_t0);
not NOT1_1782 (N6803, N5747_t0);
not NOT1_1783 (N6806, N5751_t0);
not NOT1_1784 (N6809, N5758_t0);
not NOT1_1785 (N6812, N5762_t0);
buf BUFF1_1786 (N6815, N5744_t0);
buf BUFF1_1787 (N6818, N5744_t1);
buf BUFF1_1788 (N6821, N5755_t0);
buf BUFF1_1789 (N6824, N5755_t1);
buf BUFF1_1790 (N6827, N5766_t0);
buf BUFF1_1791 (N6830, N5766_t1);
and AND4_1792 (N6833, N5850_t0, N5789_t0, N5778_t0, N5771_t0);
and AND2_1793 (N6836, N5771_t1, N3169_t0);
and AND3_1794 (N6837, N5778_t1, N5771_t2, N3173_t0);
and AND4_1795 (N6838, N5789_t1, N5771_t3, N3178_t1, N5778_t2);
and AND2_1796 (N6839, N5778_t3, N3173_t1);
and AND3_1797 (N6840, N5789_t2, N3178_t2, N5778_t4);
and AND3_1798 (N6841, N5850_t1, N5789_t3, N5778_t5);
and AND2_1799 (N6842, N5778_t6, N3173_t2);
and AND3_1800 (N6843, N5789_t4, N3178_t3, N5778_t7);
and AND2_1801 (N6844, N5789_t5, N3178_t4);
and AND5_1802 (N6845, N5856_t0, N5837_t0, N5821_t0, N5807_t0, N5799_t0);
and AND2_1803 (N6848, N5799_t1, N3185_t0);
and AND3_1804 (N6849, N5807_t1, N5799_t2, N3189_t0);
and AND4_1805 (N6850, N5821_t1, N5799_t3, N3195_t0, N5807_t2);
and AND5_1806 (N6851, N5837_t1, N5821_t2, N5799_t4, N3202_t1, N5807_t3);
and AND2_1807 (N6852, N5807_t4, N3189_t1);
and AND3_1808 (N6853, N5821_t3, N3195_t1, N5807_t5);
and AND4_1809 (N6854, N5837_t2, N5821_t4, N3202_t2, N5807_t6);
and AND4_1810 (N6855, N5856_t1, N5821_t5, N5807_t7, N5837_t3);
and AND2_1811 (N6856, N5807_t8, N3189_t2);
and AND3_1812 (N6857, N5821_t6, N3195_t2, N5807_t9);
and AND4_1813 (N6858, N5837_t4, N5821_t7, N3202_t3, N5807_t10);
and AND2_1814 (N6859, N5821_t8, N3195_t3);
and AND3_1815 (N6860, N5837_t5, N5821_t9, N3202_t4);
and AND3_1816 (N6861, N5856_t2, N5821_t10, N5837_t6);
and AND2_1817 (N6862, N5821_t11, N3195_t4);
and AND3_1818 (N6863, N5837_t7, N5821_t12, N3202_t5);
and AND2_1819 (N6864, N5837_t8, N3202_t6);
and AND2_1820 (N6865, N5850_t2, N5789_t6);
and AND2_1821 (N6866, N5856_t3, N5837_t9);
and AND4_1822 (N6867, N5870_t0, N5892_t1, N5881_t0, N5863_t0);
and AND2_1823 (N6870, N5863_t1, N3211_t0);
and AND3_1824 (N6871, N5870_t1, N5863_t2, N3215_t0);
and AND4_1825 (N6872, N5881_t1, N5863_t3, N3221_t1, N5870_t2);
and AND2_1826 (N6873, N5870_t3, N3215_t1);
and AND3_1827 (N6874, N5881_t2, N3221_t2, N5870_t4);
and AND3_1828 (N6875, N5892_t2, N5881_t3, N5870_t5);
and AND2_1829 (N6876, N5870_t6, N3215_t2);
and AND3_1830 (N6877, N3221_t3, N5881_t4, N5870_t7);
and AND2_1831 (N6878, N5881_t5, N3221_t4);
and AND2_1832 (N6879, N5892_t3, N5881_t6);
and AND2_1833 (N6880, N5881_t7, N3221_t5);
and AND5_1834 (N6881, N5905_t0, N5936_t0, N5915_t0, N5898_t0, N5926_t0);
and AND2_1835 (N6884, N5898_t1, N3229_t0);
and AND3_1836 (N6885, N5905_t1, N5898_t2, N3232_t0);
and AND4_1837 (N6886, N5915_t1, N5898_t3, N3236_t0, N5905_t2);
and AND5_1838 (N6887, N5926_t1, N5915_t2, N5898_t4, N3241_t0, N5905_t3);
and AND2_1839 (N6888, N5905_t4, N3232_t1);
and AND3_1840 (N6889, N5915_t3, N3236_t1, N5905_t5);
and AND4_1841 (N6890, N5926_t2, N5915_t4, N3241_t1, N5905_t6);
and AND2_1842 (N6891, N3236_t2, N5915_t5);
and AND3_1843 (N6892, N5926_t3, N5915_t6, N3241_t2);
and AND2_1844 (N6893, N5926_t4, N3241_t3);
nand NAND2_1845 (N6894, N5944, N6540);
nand NAND2_1846 (N6901, N5946, N6541);
nand NAND2_1847 (N6912, N5948, N6542);
nand NAND2_1848 (N6923, N5950, N6543);
nand NAND2_1849 (N6929, N5952, N6544);
nand NAND2_1850 (N6936, N5954, N6545);
nand NAND2_1851 (N6946, N5956, N6546);
nand NAND2_1852 (N6957, N5958, N6547);
nand NAND2_1853 (N6967, N6204_t0, N4575);
not NOT1_1854 (N6968, N6204_t1);
not NOT1_1855 (N6969, N6207_t0);
nand NAND2_1856 (N6970, N5967, N6555);
nand NAND2_1857 (N6977, N5969, N6556);
nand NAND2_1858 (N6988, N5971, N6557);
nand NAND2_1859 (N6998, N5973, N6558);
nand NAND2_1860 (N7006, N5975, N6559);
nand NAND2_1861 (N7020, N5977, N6560);
nand NAND2_1862 (N7036, N5979, N6561);
nand NAND2_1863 (N7049, N5989, N6569);
nand NAND2_1864 (N7055, N6210_t0, N4610);
not NOT1_1865 (N7056, N6210_t1);
and AND4_1866 (N7057, N6021, N6000_t0, N5996_t0, N5991_t0);
and AND2_1867 (N7060, N5991_t1, N3362);
and AND3_1868 (N7061, N5996_t1, N5991_t2, N3363);
and AND4_1869 (N7062, N6000_t1, N5991_t3, N3364, N5996_t2);
and AND5_1870 (N7063, N6022, N6018_t0, N6014_t0, N6009_t0, N6003_t0);
and AND2_1871 (N7064, N6003_t1, N3366);
and AND3_1872 (N7065, N6009_t1, N6003_t2, N3367);
and AND4_1873 (N7066, N6014_t1, N6003_t3, N3368, N6009_t2);
and AND5_1874 (N7067, N6018_t1, N6014_t2, N6003_t4, N3369, N6009_t3);
nand NAND2_1875 (N7068, N6594, N6024);
nand NAND2_1876 (N7073, N6595, N6026);
nand NAND2_1877 (N7077, N6596, N6028);
nand NAND2_1878 (N7080, N6597, N6030);
nand NAND2_1879 (N7086, N6598, N6599);
nand NAND2_1880 (N7091, N6600, N6601);
nand NAND2_1881 (N7095, N6602, N6603);
nand NAND2_1882 (N7098, N6604, N6038);
nand NAND2_1883 (N7099, N6605, N6606);
and AND5_1884 (N7100, N6059, N6056_t0, N6052_t0, N6047_t0, N6041_t0);
and AND2_1885 (N7103, N6041_t1, N3371);
and AND3_1886 (N7104, N6047_t1, N6041_t2, N3372);
and AND4_1887 (N7105, N6052_t1, N6041_t3, N3373, N6047_t2);
and AND5_1888 (N7106, N6056_t1, N6052_t2, N6041_t4, N3374, N6047_t3);
nand NAND2_1889 (N7107, N6060, N6621);
nand NAND2_1890 (N7114, N6062, N6622);
nand NAND2_1891 (N7125, N6064, N6623);
nand NAND2_1892 (N7136, N6066, N6624);
nand NAND2_1893 (N7142, N6068, N6625);
nand NAND2_1894 (N7149, N6070, N6626);
nand NAND2_1895 (N7159, N6072, N6627);
nand NAND2_1896 (N7170, N6074, N6628);
nand NAND2_1897 (N7180, N6076, N6629);
not NOT1_1898 (N7187, N6220_t0);
not NOT1_1899 (N7188, N6079_t0);
not NOT1_1900 (N7191, N6083_t0);
nand NAND2_1901 (N7194, N6639, N6091);
nand NAND2_1902 (N7198, N6640, N6641);
nand NAND2_1903 (N7202, N6642, N6643);
nand NAND2_1904 (N7205, N6644, N6097);
nand NAND2_1905 (N7209, N6645, N6646);
nand NAND2_1906 (N7213, N6647, N6648);
buf BUFF1_1907 (N7216, N6087_t0);
buf BUFF1_1908 (N7219, N6087_t1);
nand NAND2_1909 (N7222, N6103, N6649);
nand NAND2_1910 (N7229, N6105, N6650);
nand NAND2_1911 (N7240, N6107, N6651);
nand NAND2_1912 (N7250, N6109, N6652);
nand NAND2_1913 (N7258, N6111, N6653);
nand NAND2_1914 (N7272, N6113, N6654);
nand NAND2_1915 (N7288, N6115, N6655);
nand NAND2_1916 (N7301, N6117, N6656);
nand NAND2_1917 (N7307, N6119, N6657);
nand NAND2_1918 (N7314, N6658, N6122);
nand NAND2_1919 (N7318, N6659, N6660);
nand NAND2_1920 (N7322, N6125, N6661);
not NOT1_1921 (N7325, N6127_t0);
not NOT1_1922 (N7328, N6131_t0);
nand NAND2_1923 (N7331, N6668, N6136);
not NOT1_1924 (N7334, N6137_t0);
not NOT1_1925 (N7337, N6141_t0);
buf BUFF1_1926 (N7340, N6145_t0);
buf BUFF1_1927 (N7343, N6145_t1);
nand NAND2_1928 (N7346, N6677, N6678);
nand NAND2_1929 (N7351, N6679, N6680);
nand NAND2_1930 (N7355, N6681, N6682);
nand NAND2_1931 (N7358, N6683, N6684);
nand NAND2_1932 (N7364, N6685, N6157);
nand NAND2_1933 (N7369, N6686, N6159);
nand NAND2_1934 (N7373, N6687, N6161);
nand NAND2_1935 (N7376, N6688, N6689);
nand NAND2_1936 (N7377, N6164, N6690);
not NOT1_1937 (N7378, N6166_t0);
not NOT1_1938 (N7381, N6170_t0);
not NOT1_1939 (N7384, N6177_t0);
nand NAND2_1940 (N7387, N6702, N6703);
nand NAND2_1941 (N7391, N6704, N6705);
nand NAND2_1942 (N7394, N6706, N6186);
nand NAND2_1943 (N7398, N6707, N6708);
nand NAND2_1944 (N7402, N6709, N6710);
buf BUFF1_1945 (N7405, N6174_t0);
buf BUFF1_1946 (N7408, N6174_t1);
buf BUFF1_1947 (N7411, N5936_t1);
buf BUFF1_1948 (N7414, N5898_t5);
buf BUFF1_1949 (N7417, N5905_t7);
buf BUFF1_1950 (N7420, N5915_t7);
buf BUFF1_1951 (N7423, N5926_t5);
buf BUFF1_1952 (N7426, N5728_t1);
buf BUFF1_1953 (N7429, N5690_t5);
buf BUFF1_1954 (N7432, N5697_t7);
buf BUFF1_1955 (N7435, N5707_t7);
buf BUFF1_1956 (N7438, N5718_t5);
nand NAND2_1957 (N7441, N6192, N6711);
nand NAND2_1958 (N7444, N6194, N6712);
buf BUFF1_1959 (N7447, N5683_t4);
buf BUFF1_1960 (N7450, N5670_t10);
buf BUFF1_1961 (N7453, N5632_t5);
buf BUFF1_1962 (N7456, N5654_t13);
buf BUFF1_1963 (N7459, N5640_t11);
buf BUFF1_1964 (N7462, N5640_t12);
buf BUFF1_1965 (N7465, N5683_t5);
buf BUFF1_1966 (N7468, N5670_t11);
buf BUFF1_1967 (N7471, N5632_t6);
buf BUFF1_1968 (N7474, N5654_t14);
not NOT1_1969 (N7477, N6196_t0);
not NOT1_1970 (N7478, N6199_t0);
buf BUFF1_1971 (N7479, N5850_t3);
buf BUFF1_1972 (N7482, N5789_t7);
buf BUFF1_1973 (N7485, N5771_t4);
buf BUFF1_1974 (N7488, N5778_t8);
buf BUFF1_1975 (N7491, N5850_t4);
buf BUFF1_1976 (N7494, N5789_t8);
buf BUFF1_1977 (N7497, N5771_t5);
buf BUFF1_1978 (N7500, N5778_t9);
buf BUFF1_1979 (N7503, N5856_t4);
buf BUFF1_1980 (N7506, N5837_t10);
buf BUFF1_1981 (N7509, N5799_t5);
buf BUFF1_1982 (N7512, N5821_t13);
buf BUFF1_1983 (N7515, N5807_t11);
buf BUFF1_1984 (N7518, N5807_t12);
buf BUFF1_1985 (N7521, N5856_t5);
buf BUFF1_1986 (N7524, N5837_t11);
buf BUFF1_1987 (N7527, N5799_t6);
buf BUFF1_1988 (N7530, N5821_t14);
buf BUFF1_1989 (N7533, N5863_t4);
buf BUFF1_1990 (N7536, N5863_t5);
buf BUFF1_1991 (N7539, N5870_t8);
buf BUFF1_1992 (N7542, N5870_t9);
buf BUFF1_1993 (N7545, N5881_t8);
buf BUFF1_1994 (N7548, N5881_t9);
not NOT1_1995 (N7551, N6214_t0);
not NOT1_1996 (N7552, N6217_t0);
buf BUFF1_1997 (N7553, N5981_t0);
not NOT1_1998 (N7556, N6249_t0);
not NOT1_1999 (N7557, N6252_t0);
not NOT1_2000 (N7558, N6243_t0);
not NOT1_2001 (N7559, N6246_t0);
nand NAND2_2002 (N7560, N6731, N6732);
nand NAND2_2003 (N7563, N6729, N6730);
nand NAND2_2004 (N7566, N6735, N6736);
nand NAND2_2005 (N7569, N6733, N6734);
not NOT1_2006 (N7572, N6232_t0);
not NOT1_2007 (N7573, N6236_t0);
nand NAND2_2008 (N7574, N6743, N6744);
nand NAND2_2009 (N7577, N6741, N6742);
not NOT1_2010 (N7580, N6263_t0);
not NOT1_2011 (N7581, N6266_t0);
nand NAND2_2012 (N7582, N6753, N6754);
nand NAND2_2013 (N7585, N6751, N6752);
nand NAND2_2014 (N7588, N6757, N6758);
nand NAND2_2015 (N7591, N6755, N6756);
or OR5_2016 (N7609, N3096, N6766, N6767, N6768, N6769);
or OR2_2017 (N7613, N3107_t5, N6782);
or OR5_2018 (N7620, N3136, N6787, N6788, N6789, N6790);
or OR4_2019 (N7649, N3168, N6836, N6837, N6838);
or OR2_2020 (N7650, N3173_t3, N6844);
or OR5_2021 (N7655, N3184, N6848, N6849, N6850, N6851);
or OR2_2022 (N7659, N3195_t5, N6864);
or OR4_2023 (N7668, N3210, N6870, N6871, N6872);
or OR5_2024 (N7671, N3228, N6884, N6885, N6886, N6887);
nand NAND2_2025 (N7744, N3661_t1, N6968);
nand NAND2_2026 (N7822, N3664_t1, N7056);
or OR4_2027 (N7825, N3361, N7060, N7061, N7062);
or OR5_2028 (N7826, N3365, N7064, N7065, N7066, N7067);
or OR5_2029 (N7852, N3370, N7103, N7104, N7105, N7106);
or OR4_2030 (N8114, N3101_t3, N6777, N6778, N6779);
or OR5_2031 (N8117, N3097_t1, N6770, N6771, N6772, N6773);
nor NOR3_2032 (N8131, N3101_t4, N6780, N6781);
nor NOR4_2033 (N8134, N3097_t2, N6774, N6775, N6776);
nand NAND2_2034 (N8144, N6199_t1, N7477);
nand NAND2_2035 (N8145, N6196_t1, N7478);
or OR4_2036 (N8146, N3169_t1, N6839, N6840, N6841);
nor NOR3_2037 (N8156, N3169_t2, N6842, N6843);
or OR4_2038 (N8166, N3189_t3, N6859, N6860, N6861);
or OR5_2039 (N8169, N3185_t1, N6852, N6853, N6854, N6855);
nor NOR3_2040 (N8183, N3189_t4, N6862, N6863);
nor NOR4_2041 (N8186, N3185_t2, N6856, N6857, N6858);
or OR4_2042 (N8196, N3211_t1, N6873, N6874, N6875);
nor NOR3_2043 (N8200, N3211_t2, N6876, N6877);
or OR3_2044 (N8204, N3215_t3, N6878, N6879);
nor NOR2_2045 (N8208, N3215_t4, N6880);
nand NAND2_2046 (N8216, N6252_t1, N7556);
nand NAND2_2047 (N8217, N6249_t1, N7557);
nand NAND2_2048 (N8218, N6246_t1, N7558);
nand NAND2_2049 (N8219, N6243_t1, N7559);
nand NAND2_2050 (N8232, N6266_t1, N7580);
nand NAND2_2051 (N8233, N6263_t1, N7581);
not NOT1_2052 (N8242, N7411_t0);
not NOT1_2053 (N8243, N7414_t0);
not NOT1_2054 (N8244, N7417_t0);
not NOT1_2055 (N8245, N7420_t0);
not NOT1_2056 (N8246, N7423_t0);
not NOT1_2057 (N8247, N7426_t0);
not NOT1_2058 (N8248, N7429_t0);
not NOT1_2059 (N8249, N7432_t0);
not NOT1_2060 (N8250, N7435_t0);
not NOT1_2061 (N8251, N7438_t0);
not NOT1_2062 (N8252, N7136_t0);
not NOT1_2063 (N8253, N6923_t0);
not NOT1_2064 (N8254, N6762_t0);
not NOT1_2065 (N8260, N7459_t0);
not NOT1_2066 (N8261, N7462_t0);
and AND2_2067 (N8262, N3122_t1, N6762_t1);
and AND2_2068 (N8269, N3155_t1, N6784_t0);
not NOT1_2069 (N8274, N6815_t0);
not NOT1_2070 (N8275, N6818_t0);
not NOT1_2071 (N8276, N6821_t0);
not NOT1_2072 (N8277, N6824_t0);
not NOT1_2073 (N8278, N6827_t0);
not NOT1_2074 (N8279, N6830_t0);
and AND3_2075 (N8280, N5740_t1, N5736_t1, N6815_t1);
and AND3_2076 (N8281, N6800_t0, N6797_t0, N6818_t1);
and AND3_2077 (N8282, N5751_t1, N5747_t1, N6821_t1);
and AND3_2078 (N8283, N6806_t0, N6803_t0, N6824_t1);
and AND3_2079 (N8284, N5762_t1, N5758_t1, N6827_t1);
and AND3_2080 (N8285, N6812_t0, N6809_t0, N6830_t1);
not NOT1_2081 (N8288, N6845_t0);
not NOT1_2082 (N8294, N7488_t0);
not NOT1_2083 (N8295, N7500_t0);
not NOT1_2084 (N8296, N7515_t0);
not NOT1_2085 (N8297, N7518_t0);
and AND2_2086 (N8298, N6833_t0, N6845_t1);
and AND2_2087 (N8307, N6867_t0, N6881_t0);
not NOT1_2088 (N8315, N7533_t0);
not NOT1_2089 (N8317, N7536_t0);
not NOT1_2090 (N8319, N7539_t0);
not NOT1_2091 (N8321, N7542_t0);
nand NAND2_2092 (N8322, N7545_t0, N4543);
not NOT1_2093 (N8323, N7545_t1);
nand NAND2_2094 (N8324, N7548_t0, N5943);
not NOT1_2095 (N8325, N7548_t1);
nand NAND2_2096 (N8326, N6967, N7744);
and AND4_2097 (N8333, N6901_t0, N6923_t1, N6912_t0, N6894_t0);
and AND2_2098 (N8337, N6894_t1, N4545_t0);
and AND3_2099 (N8338, N6901_t1, N6894_t2, N4549_t0);
and AND4_2100 (N8339, N6912_t1, N6894_t3, N4555_t1, N6901_t2);
and AND2_2101 (N8340, N6901_t3, N4549_t1);
and AND3_2102 (N8341, N6912_t2, N4555_t2, N6901_t4);
and AND3_2103 (N8342, N6923_t2, N6912_t3, N6901_t5);
and AND2_2104 (N8343, N6901_t6, N4549_t2);
and AND3_2105 (N8344, N4555_t3, N6912_t4, N6901_t7);
and AND2_2106 (N8345, N6912_t5, N4555_t4);
and AND2_2107 (N8346, N6923_t3, N6912_t6);
and AND2_2108 (N8347, N6912_t7, N4555_t5);
and AND2_2109 (N8348, N6929_t0, N4563_t0);
and AND3_2110 (N8349, N6936_t0, N6929_t1, N4566_t0);
and AND4_2111 (N8350, N6946_t0, N6929_t2, N4570_t0, N6936_t1);
and AND5_2112 (N8351, N6957_t0, N6946_t1, N6929_t3, N5960_t0, N6936_t2);
and AND2_2113 (N8352, N6936_t3, N4566_t1);
and AND3_2114 (N8353, N6946_t2, N4570_t1, N6936_t4);
and AND4_2115 (N8354, N6957_t1, N6946_t3, N5960_t1, N6936_t5);
and AND2_2116 (N8355, N4570_t2, N6946_t4);
and AND3_2117 (N8356, N6957_t2, N6946_t5, N5960_t2);
and AND2_2118 (N8357, N6957_t3, N5960_t3);
nand NAND2_2119 (N8358, N7055, N7822);
and AND4_2120 (N8365, N7049_t0, N6988_t0, N6977_t0, N6970_t0);
and AND2_2121 (N8369, N6970_t1, N4577_t0);
and AND3_2122 (N8370, N6977_t1, N6970_t2, N4581_t0);
and AND4_2123 (N8371, N6988_t1, N6970_t3, N4586_t1, N6977_t2);
and AND2_2124 (N8372, N6977_t3, N4581_t1);
and AND3_2125 (N8373, N6988_t2, N4586_t2, N6977_t4);
and AND3_2126 (N8374, N7049_t1, N6988_t3, N6977_t5);
and AND2_2127 (N8375, N6977_t6, N4581_t2);
and AND3_2128 (N8376, N6988_t4, N4586_t3, N6977_t7);
and AND2_2129 (N8377, N6988_t5, N4586_t4);
and AND2_2130 (N8378, N6998_t0, N4593_t0);
and AND3_2131 (N8379, N7006_t0, N6998_t1, N4597_t0);
and AND4_2132 (N8380, N7020_t0, N6998_t2, N4603_t0, N7006_t1);
and AND5_2133 (N8381, N7036_t0, N7020_t1, N6998_t3, N5981_t1, N7006_t2);
and AND2_2134 (N8382, N7006_t3, N4597_t1);
and AND3_2135 (N8383, N7020_t2, N4603_t1, N7006_t4);
and AND4_2136 (N8384, N7036_t1, N7020_t3, N5981_t2, N7006_t5);
and AND2_2137 (N8385, N7006_t6, N4597_t2);
and AND3_2138 (N8386, N7020_t4, N4603_t2, N7006_t7);
and AND4_2139 (N8387, N7036_t2, N7020_t5, N5981_t3, N7006_t8);
and AND2_2140 (N8388, N7020_t6, N4603_t3);
and AND3_2141 (N8389, N7036_t3, N7020_t7, N5981_t4);
and AND2_2142 (N8390, N7020_t8, N4603_t4);
and AND3_2143 (N8391, N7036_t4, N7020_t9, N5981_t5);
and AND2_2144 (N8392, N7036_t5, N5981_t6);
and AND2_2145 (N8393, N7049_t2, N6988_t6);
and AND2_2146 (N8394, N7057_t0, N7063);
and AND2_2147 (N8404, N7057_t1, N7826);
and AND4_2148 (N8405, N7098, N7077_t0, N7073_t0, N7068_t0);
and AND2_2149 (N8409, N7068_t1, N4632);
and AND3_2150 (N8410, N7073_t1, N7068_t2, N4634);
and AND4_2151 (N8411, N7077_t1, N7068_t3, N4635, N7073_t2);
and AND5_2152 (N8412, N7099, N7095_t0, N7091_t0, N7086_t0, N7080_t0);
and AND2_2153 (N8415, N7080_t1, N4638);
and AND3_2154 (N8416, N7086_t1, N7080_t2, N4639);
and AND4_2155 (N8417, N7091_t1, N7080_t3, N4640, N7086_t2);
and AND5_2156 (N8418, N7095_t1, N7091_t2, N7080_t4, N4641, N7086_t3);
and AND2_2157 (N8421, N3375_t1, N7100_t0);
and AND4_2158 (N8430, N7114_t0, N7136_t1, N7125_t0, N7107_t0);
and AND2_2159 (N8433, N7107_t1, N4657_t0);
and AND3_2160 (N8434, N7114_t1, N7107_t2, N4661_t0);
and AND4_2161 (N8435, N7125_t1, N7107_t3, N4667_t1, N7114_t2);
and AND2_2162 (N8436, N7114_t3, N4661_t1);
and AND3_2163 (N8437, N7125_t2, N4667_t2, N7114_t4);
and AND3_2164 (N8438, N7136_t2, N7125_t3, N7114_t5);
and AND2_2165 (N8439, N7114_t6, N4661_t2);
and AND3_2166 (N8440, N4667_t3, N7125_t4, N7114_t7);
and AND2_2167 (N8441, N7125_t5, N4667_t4);
and AND2_2168 (N8442, N7136_t3, N7125_t6);
and AND2_2169 (N8443, N7125_t7, N4667_t5);
and AND5_2170 (N8444, N7149_t0, N7180_t0, N7159_t0, N7142_t0, N7170_t0);
and AND2_2171 (N8447, N7142_t1, N4675_t0);
and AND3_2172 (N8448, N7149_t1, N7142_t2, N4678_t0);
and AND4_2173 (N8449, N7159_t1, N7142_t3, N4682_t0, N7149_t2);
and AND5_2174 (N8450, N7170_t1, N7159_t2, N7142_t4, N4687_t0, N7149_t3);
and AND2_2175 (N8451, N7149_t4, N4678_t1);
and AND3_2176 (N8452, N7159_t3, N4682_t1, N7149_t5);
and AND4_2177 (N8453, N7170_t2, N7159_t4, N4687_t1, N7149_t6);
and AND2_2178 (N8454, N4682_t2, N7159_t5);
and AND3_2179 (N8455, N7170_t3, N7159_t6, N4687_t2);
and AND2_2180 (N8456, N7170_t4, N4687_t3);
not NOT1_2181 (N8457, N7194_t0);
not NOT1_2182 (N8460, N7198_t0);
not NOT1_2183 (N8463, N7205_t0);
not NOT1_2184 (N8466, N7209_t0);
not NOT1_2185 (N8469, N7216_t0);
not NOT1_2186 (N8470, N7219_t0);
buf BUFF1_2187 (N8471, N7202_t0);
buf BUFF1_2188 (N8474, N7202_t1);
buf BUFF1_2189 (N8477, N7213_t0);
buf BUFF1_2190 (N8480, N7213_t1);
and AND3_2191 (N8483, N6083_t1, N6079_t1, N7216_t1);
and AND3_2192 (N8484, N7191_t0, N7188_t0, N7219_t1);
and AND4_2193 (N8485, N7301_t0, N7240_t0, N7229_t0, N7222_t0);
and AND2_2194 (N8488, N7222_t1, N4702_t0);
and AND3_2195 (N8489, N7229_t1, N7222_t2, N4706_t0);
and AND4_2196 (N8490, N7240_t1, N7222_t3, N4711_t1, N7229_t2);
and AND2_2197 (N8491, N7229_t3, N4706_t1);
and AND3_2198 (N8492, N7240_t2, N4711_t2, N7229_t4);
and AND3_2199 (N8493, N7301_t1, N7240_t3, N7229_t5);
and AND2_2200 (N8494, N7229_t6, N4706_t2);
and AND3_2201 (N8495, N7240_t4, N4711_t3, N7229_t7);
and AND2_2202 (N8496, N7240_t5, N4711_t4);
and AND5_2203 (N8497, N7307_t0, N7288_t0, N7272_t0, N7258_t0, N7250_t0);
and AND2_2204 (N8500, N7250_t1, N4718_t0);
and AND3_2205 (N8501, N7258_t1, N7250_t2, N4722_t0);
and AND4_2206 (N8502, N7272_t1, N7250_t3, N4728_t0, N7258_t2);
and AND5_2207 (N8503, N7288_t1, N7272_t2, N7250_t4, N4735_t1, N7258_t3);
and AND2_2208 (N8504, N7258_t4, N4722_t1);
and AND3_2209 (N8505, N7272_t3, N4728_t1, N7258_t5);
and AND4_2210 (N8506, N7288_t2, N7272_t4, N4735_t2, N7258_t6);
and AND4_2211 (N8507, N7307_t1, N7272_t5, N7258_t7, N7288_t3);
and AND2_2212 (N8508, N7258_t8, N4722_t2);
and AND3_2213 (N8509, N7272_t6, N4728_t2, N7258_t9);
and AND4_2214 (N8510, N7288_t4, N7272_t7, N4735_t3, N7258_t10);
and AND2_2215 (N8511, N7272_t8, N4728_t3);
and AND3_2216 (N8512, N7288_t5, N7272_t9, N4735_t4);
and AND3_2217 (N8513, N7307_t2, N7272_t10, N7288_t6);
and AND2_2218 (N8514, N7272_t11, N4728_t4);
and AND3_2219 (N8515, N7288_t7, N7272_t12, N4735_t5);
and AND2_2220 (N8516, N7288_t8, N4735_t6);
and AND2_2221 (N8517, N7301_t2, N7240_t6);
and AND2_2222 (N8518, N7307_t3, N7288_t9);
not NOT1_2223 (N8519, N7314_t0);
not NOT1_2224 (N8522, N7318_t0);
buf BUFF1_2225 (N8525, N7322_t0);
buf BUFF1_2226 (N8528, N7322_t1);
buf BUFF1_2227 (N8531, N7331_t0);
buf BUFF1_2228 (N8534, N7331_t1);
not NOT1_2229 (N8537, N7340_t0);
not NOT1_2230 (N8538, N7343_t0);
and AND3_2231 (N8539, N6141_t1, N6137_t1, N7340_t1);
and AND3_2232 (N8540, N7337_t0, N7334_t0, N7343_t1);
and AND4_2233 (N8541, N7376, N7355_t0, N7351_t0, N7346_t0);
and AND2_2234 (N8545, N7346_t1, N4757);
and AND3_2235 (N8546, N7351_t1, N7346_t2, N4758);
and AND4_2236 (N8547, N7355_t1, N7346_t3, N4759, N7351_t2);
and AND5_2237 (N8548, N7377, N7373_t0, N7369_t0, N7364_t0, N7358_t0);
and AND2_2238 (N8551, N7358_t1, N4762);
and AND3_2239 (N8552, N7364_t1, N7358_t2, N4764);
and AND4_2240 (N8553, N7369_t1, N7358_t3, N4766, N7364_t2);
and AND5_2241 (N8554, N7373_t1, N7369_t2, N7358_t4, N4767, N7364_t3);
not NOT1_2242 (N8555, N7387_t0);
not NOT1_2243 (N8558, N7394_t0);
not NOT1_2244 (N8561, N7398_t0);
not NOT1_2245 (N8564, N7405_t0);
not NOT1_2246 (N8565, N7408_t0);
buf BUFF1_2247 (N8566, N7391_t0);
buf BUFF1_2248 (N8569, N7391_t1);
buf BUFF1_2249 (N8572, N7402_t0);
buf BUFF1_2250 (N8575, N7402_t1);
and AND3_2251 (N8578, N6170_t1, N6166_t1, N7405_t1);
and AND3_2252 (N8579, N7381_t0, N7378_t0, N7408_t1);
buf BUFF1_2253 (N8580, N7180_t1);
buf BUFF1_2254 (N8583, N7142_t5);
buf BUFF1_2255 (N8586, N7149_t7);
buf BUFF1_2256 (N8589, N7159_t7);
buf BUFF1_2257 (N8592, N7170_t5);
buf BUFF1_2258 (N8595, N6929_t4);
buf BUFF1_2259 (N8598, N6936_t6);
buf BUFF1_2260 (N8601, N6946_t6);
buf BUFF1_2261 (N8604, N6957_t4);
not NOT1_2262 (N8607, N7441_t0);
nand NAND2_2263 (N8608, N7441_t1, N5469);
not NOT1_2264 (N8609, N7444_t0);
nand NAND2_2265 (N8610, N7444_t1, N4793);
not NOT1_2266 (N8615, N7447_t0);
not NOT1_2267 (N8616, N7450_t0);
not NOT1_2268 (N8617, N7453_t0);
not NOT1_2269 (N8618, N7456_t0);
not NOT1_2270 (N8619, N7474_t0);
not NOT1_2271 (N8624, N7465_t0);
not NOT1_2272 (N8625, N7468_t0);
not NOT1_2273 (N8626, N7471_t0);
nand NAND2_2274 (N8627, N8144, N8145);
not NOT1_2275 (N8632, N7479_t0);
not NOT1_2276 (N8633, N7482_t0);
not NOT1_2277 (N8634, N7485_t0);
not NOT1_2278 (N8637, N7491_t0);
not NOT1_2279 (N8638, N7494_t0);
not NOT1_2280 (N8639, N7497_t0);
not NOT1_2281 (N8644, N7503_t0);
not NOT1_2282 (N8645, N7506_t0);
not NOT1_2283 (N8646, N7509_t0);
not NOT1_2284 (N8647, N7512_t0);
not NOT1_2285 (N8648, N7530_t0);
not NOT1_2286 (N8653, N7521_t0);
not NOT1_2287 (N8654, N7524_t0);
not NOT1_2288 (N8655, N7527_t0);
buf BUFF1_2289 (N8660, N6894_t4);
buf BUFF1_2290 (N8663, N6894_t5);
buf BUFF1_2291 (N8666, N6901_t8);
buf BUFF1_2292 (N8669, N6901_t9);
buf BUFF1_2293 (N8672, N6912_t8);
buf BUFF1_2294 (N8675, N6912_t9);
buf BUFF1_2295 (N8678, N7049_t3);
buf BUFF1_2296 (N8681, N6988_t7);
buf BUFF1_2297 (N8684, N6970_t4);
buf BUFF1_2298 (N8687, N6977_t8);
buf BUFF1_2299 (N8690, N7049_t4);
buf BUFF1_2300 (N8693, N6988_t8);
buf BUFF1_2301 (N8696, N6970_t5);
buf BUFF1_2302 (N8699, N6977_t9);
buf BUFF1_2303 (N8702, N7036_t6);
buf BUFF1_2304 (N8705, N6998_t4);
buf BUFF1_2305 (N8708, N7020_t10);
buf BUFF1_2306 (N8711, N7006_t9);
buf BUFF1_2307 (N8714, N7006_t10);
not NOT1_2308 (N8717, N7553_t0);
buf BUFF1_2309 (N8718, N7036_t7);
buf BUFF1_2310 (N8721, N6998_t5);
buf BUFF1_2311 (N8724, N7020_t11);
nand NAND2_2312 (N8727, N8216, N8217);
nand NAND2_2313 (N8730, N8218, N8219);
not NOT1_2314 (N8733, N7574_t0);
not NOT1_2315 (N8734, N7577_t0);
buf BUFF1_2316 (N8735, N7107_t4);
buf BUFF1_2317 (N8738, N7107_t5);
buf BUFF1_2318 (N8741, N7114_t8);
buf BUFF1_2319 (N8744, N7114_t9);
buf BUFF1_2320 (N8747, N7125_t8);
buf BUFF1_2321 (N8750, N7125_t9);
not NOT1_2322 (N8753, N7560_t0);
not NOT1_2323 (N8754, N7563_t0);
not NOT1_2324 (N8755, N7566_t0);
not NOT1_2325 (N8756, N7569_t0);
buf BUFF1_2326 (N8757, N7301_t3);
buf BUFF1_2327 (N8760, N7240_t7);
buf BUFF1_2328 (N8763, N7222_t4);
buf BUFF1_2329 (N8766, N7229_t8);
buf BUFF1_2330 (N8769, N7301_t4);
buf BUFF1_2331 (N8772, N7240_t8);
buf BUFF1_2332 (N8775, N7222_t5);
buf BUFF1_2333 (N8778, N7229_t9);
buf BUFF1_2334 (N8781, N7307_t4);
buf BUFF1_2335 (N8784, N7288_t10);
buf BUFF1_2336 (N8787, N7250_t5);
buf BUFF1_2337 (N8790, N7272_t13);
buf BUFF1_2338 (N8793, N7258_t11);
buf BUFF1_2339 (N8796, N7258_t12);
buf BUFF1_2340 (N8799, N7307_t5);
buf BUFF1_2341 (N8802, N7288_t11);
buf BUFF1_2342 (N8805, N7250_t6);
buf BUFF1_2343 (N8808, N7272_t14);
nand NAND2_2344 (N8811, N8232, N8233);
not NOT1_2345 (N8814, N7588_t0);
not NOT1_2346 (N8815, N7591_t0);
not NOT1_2347 (N8816, N7582_t0);
not NOT1_2348 (N8817, N7585_t0);
and AND2_2349 (N8818, N7620_t0, N3155_t2);
and AND2_2350 (N8840, N3122_t2, N7609_t0);
not NOT1_2351 (N8857, N7609_t1);
and AND3_2352 (N8861, N6797_t1, N5740_t2, N8274);
and AND3_2353 (N8862, N5736_t2, N6800_t1, N8275);
and AND3_2354 (N8863, N6803_t1, N5751_t2, N8276);
and AND3_2355 (N8864, N5747_t2, N6806_t1, N8277);
and AND3_2356 (N8865, N6809_t1, N5762_t2, N8278);
and AND3_2357 (N8866, N5758_t2, N6812_t1, N8279);
not NOT1_2358 (N8871, N7655_t0);
and AND2_2359 (N8874, N6833_t1, N7655_t1);
and AND2_2360 (N8878, N7671_t0, N6867_t1);
not NOT1_2361 (N8879, N8196_t0);
nand NAND2_2362 (N8880, N8196_t1, N8315);
not NOT1_2363 (N8881, N8200_t0);
nand NAND2_2364 (N8882, N8200_t1, N8317);
not NOT1_2365 (N8883, N8204_t0);
nand NAND2_2366 (N8884, N8204_t1, N8319);
not NOT1_2367 (N8885, N8208_t0);
nand NAND2_2368 (N8886, N8208_t1, N8321);
nand NAND2_2369 (N8887, N3658_t1, N8323);
nand NAND2_2370 (N8888, N4817_t1, N8325);
or OR4_2371 (N8898, N4544, N8337, N8338, N8339);
or OR5_2372 (N8902, N4562, N8348, N8349, N8350, N8351);
or OR4_2373 (N8920, N4576, N8369, N8370, N8371);
or OR2_2374 (N8924, N4581_t3, N8377);
or OR5_2375 (N8927, N4592, N8378, N8379, N8380, N8381);
or OR2_2376 (N8931, N4603_t5, N8392);
or OR2_2377 (N8943, N7825, N8404);
or OR4_2378 (N8950, N4630, N8409, N8410, N8411);
or OR5_2379 (N8956, N4637, N8415, N8416, N8417, N8418);
not NOT1_2380 (N8959, N7852_t0);
and AND2_2381 (N8960, N3375_t2, N7852_t1);
or OR4_2382 (N8963, N4656, N8433, N8434, N8435);
or OR5_2383 (N8966, N4674, N8447, N8448, N8449, N8450);
and AND3_2384 (N8991, N7188_t1, N6083_t2, N8469);
and AND3_2385 (N8992, N6079_t2, N7191_t1, N8470);
or OR4_2386 (N8995, N4701, N8488, N8489, N8490);
or OR2_2387 (N8996, N4706_t3, N8496);
or OR5_2388 (N9001, N4717, N8500, N8501, N8502, N8503);
or OR2_2389 (N9005, N4728_t5, N8516);
and AND3_2390 (N9024, N7334_t1, N6141_t2, N8537);
and AND3_2391 (N9025, N6137_t2, N7337_t1, N8538);
or OR4_2392 (N9029, N4756, N8545, N8546, N8547);
or OR5_2393 (N9035, N4760, N8551, N8552, N8553, N8554);
and AND3_2394 (N9053, N7378_t1, N6170_t2, N8564);
and AND3_2395 (N9054, N6166_t2, N7381_t1, N8565);
nand NAND2_2396 (N9064, N4303_t1, N8607);
nand NAND2_2397 (N9065, N3507_t1, N8609);
not NOT1_2398 (N9066, N8114_t0);
nand NAND2_2399 (N9067, N8114_t1, N4795);
or OR2_2400 (N9068, N7613_t0, N6783);
not NOT1_2401 (N9071, N8117_t0);
not NOT1_2402 (N9072, N8131_t0);
nand NAND2_2403 (N9073, N8131_t1, N6195);
not NOT1_2404 (N9074, N7613_t1);
not NOT1_2405 (N9077, N8134_t0);
or OR2_2406 (N9079, N7650_t0, N6865);
not NOT1_2407 (N9082, N8146_t0);
not NOT1_2408 (N9083, N7650_t1);
not NOT1_2409 (N9086, N8156_t0);
not NOT1_2410 (N9087, N8166_t0);
nand NAND2_2411 (N9088, N8166_t1, N4813);
or OR2_2412 (N9089, N7659_t0, N6866);
not NOT1_2413 (N9092, N8169_t0);
not NOT1_2414 (N9093, N8183_t0);
nand NAND2_2415 (N9094, N8183_t1, N6203);
not NOT1_2416 (N9095, N7659_t1);
not NOT1_2417 (N9098, N8186_t0);
or OR4_2418 (N9099, N4545_t1, N8340, N8341, N8342);
nor NOR3_2419 (N9103, N4545_t2, N8343, N8344);
or OR3_2420 (N9107, N4549_t3, N8345, N8346);
nor NOR2_2421 (N9111, N4549_t4, N8347);
or OR4_2422 (N9117, N4577_t1, N8372, N8373, N8374);
nor NOR3_2423 (N9127, N4577_t2, N8375, N8376);
nor NOR3_2424 (N9146, N4597_t3, N8390, N8391);
nor NOR4_2425 (N9149, N4593_t1, N8385, N8386, N8387);
nand NAND2_2426 (N9159, N7577_t1, N8733);
nand NAND2_2427 (N9160, N7574_t1, N8734);
or OR4_2428 (N9161, N4657_t1, N8436, N8437, N8438);
nor NOR3_2429 (N9165, N4657_t2, N8439, N8440);
or OR3_2430 (N9169, N4661_t3, N8441, N8442);
nor NOR2_2431 (N9173, N4661_t4, N8443);
nand NAND2_2432 (N9179, N7563_t1, N8753);
nand NAND2_2433 (N9180, N7560_t1, N8754);
nand NAND2_2434 (N9181, N7569_t1, N8755);
nand NAND2_2435 (N9182, N7566_t1, N8756);
or OR4_2436 (N9183, N4702_t1, N8491, N8492, N8493);
nor NOR3_2437 (N9193, N4702_t2, N8494, N8495);
or OR4_2438 (N9203, N4722_t3, N8511, N8512, N8513);
or OR5_2439 (N9206, N4718_t1, N8504, N8505, N8506, N8507);
nor NOR3_2440 (N9220, N4722_t4, N8514, N8515);
nor NOR4_2441 (N9223, N4718_t2, N8508, N8509, N8510);
nand NAND2_2442 (N9234, N7591_t1, N8814);
nand NAND2_2443 (N9235, N7588_t1, N8815);
nand NAND2_2444 (N9236, N7585_t1, N8816);
nand NAND2_2445 (N9237, N7582_t1, N8817);
or OR2_2446 (N9238, N3159_t1, N8818);
or OR2_2447 (N9242, N3126_t1, N8840);
nand NAND2_2448 (N9243, N8324, N8888);
not NOT1_2449 (N9244, N8580_t0);
not NOT1_2450 (N9245, N8583_t0);
not NOT1_2451 (N9246, N8586_t0);
not NOT1_2452 (N9247, N8589_t0);
not NOT1_2453 (N9248, N8592_t0);
not NOT1_2454 (N9249, N8595_t0);
not NOT1_2455 (N9250, N8598_t0);
not NOT1_2456 (N9251, N8601_t0);
not NOT1_2457 (N9252, N8604_t0);
nor NOR2_2458 (N9256, N8861, N8280);
nor NOR2_2459 (N9257, N8862, N8281);
nor NOR2_2460 (N9258, N8863, N8282);
nor NOR2_2461 (N9259, N8864, N8283);
nor NOR2_2462 (N9260, N8865, N8284);
nor NOR2_2463 (N9261, N8866, N8285);
not NOT1_2464 (N9262, N8627_t0);
or OR2_2465 (N9265, N7649, N8874);
or OR2_2466 (N9268, N7668, N8878);
nand NAND2_2467 (N9271, N7533_t1, N8879);
nand NAND2_2468 (N9272, N7536_t1, N8881);
nand NAND2_2469 (N9273, N7539_t1, N8883);
nand NAND2_2470 (N9274, N7542_t1, N8885);
nand NAND2_2471 (N9275, N8322, N8887);
not NOT1_2472 (N9276, N8333_t0);
and AND5_2473 (N9280, N6936_t7, N8326_t0, N6946_t7, N6929_t5, N6957_t5);
and AND5_2474 (N9285, N367_t2, N8326_t1, N6946_t8, N6957_t6, N6936_t8);
and AND4_2475 (N9286, N367_t3, N8326_t2, N6946_t9, N6957_t7);
and AND3_2476 (N9287, N367_t4, N8326_t3, N6957_t8);
and AND2_2477 (N9288, N367_t5, N8326_t4);
not NOT1_2478 (N9290, N8660_t0);
not NOT1_2479 (N9292, N8663_t0);
not NOT1_2480 (N9294, N8666_t0);
not NOT1_2481 (N9296, N8669_t0);
nand NAND2_2482 (N9297, N8672_t0, N5966);
not NOT1_2483 (N9298, N8672_t1);
nand NAND2_2484 (N9299, N8675_t0, N6969);
not NOT1_2485 (N9300, N8675_t1);
not NOT1_2486 (N9301, N8365_t0);
and AND5_2487 (N9307, N8358_t0, N7036_t8, N7020_t12, N7006_t11, N6998_t6);
and AND4_2488 (N9314, N8358_t1, N7020_t13, N7006_t12, N7036_t9);
and AND3_2489 (N9315, N8358_t2, N7020_t14, N7036_t10);
and AND2_2490 (N9318, N8358_t3, N7036_t11);
not NOT1_2491 (N9319, N8687_t0);
not NOT1_2492 (N9320, N8699_t0);
not NOT1_2493 (N9321, N8711_t0);
not NOT1_2494 (N9322, N8714_t0);
not NOT1_2495 (N9323, N8727_t0);
not NOT1_2496 (N9324, N8730_t0);
not NOT1_2497 (N9326, N8405_t0);
and AND2_2498 (N9332, N8405_t1, N8412_t0);
or OR2_2499 (N9339, N4193_t1, N8960);
and AND2_2500 (N9344, N8430_t0, N8444_t0);
not NOT1_2501 (N9352, N8735_t0);
not NOT1_2502 (N9354, N8738_t0);
not NOT1_2503 (N9356, N8741_t0);
not NOT1_2504 (N9358, N8744_t0);
nand NAND2_2505 (N9359, N8747_t0, N6078);
not NOT1_2506 (N9360, N8747_t1);
nand NAND2_2507 (N9361, N8750_t0, N7187);
not NOT1_2508 (N9362, N8750_t1);
not NOT1_2509 (N9363, N8471_t0);
not NOT1_2510 (N9364, N8474_t0);
not NOT1_2511 (N9365, N8477_t0);
not NOT1_2512 (N9366, N8480_t0);
nor NOR2_2513 (N9367, N8991, N8483);
nor NOR2_2514 (N9368, N8992, N8484);
and AND3_2515 (N9369, N7198_t1, N7194_t1, N8471_t1);
and AND3_2516 (N9370, N8460_t0, N8457_t0, N8474_t1);
and AND3_2517 (N9371, N7209_t1, N7205_t1, N8477_t1);
and AND3_2518 (N9372, N8466_t0, N8463_t0, N8480_t1);
not NOT1_2519 (N9375, N8497_t0);
not NOT1_2520 (N9381, N8766_t0);
not NOT1_2521 (N9382, N8778_t0);
not NOT1_2522 (N9383, N8793_t0);
not NOT1_2523 (N9384, N8796_t0);
and AND2_2524 (N9385, N8485_t0, N8497_t1);
not NOT1_2525 (N9392, N8525_t0);
not NOT1_2526 (N9393, N8528_t0);
not NOT1_2527 (N9394, N8531_t0);
not NOT1_2528 (N9395, N8534_t0);
and AND3_2529 (N9396, N7318_t1, N7314_t1, N8525_t1);
and AND3_2530 (N9397, N8522_t0, N8519_t0, N8528_t1);
and AND3_2531 (N9398, N6131_t1, N6127_t1, N8531_t1);
and AND3_2532 (N9399, N7328_t0, N7325_t0, N8534_t1);
nor NOR2_2533 (N9400, N9024, N8539);
nor NOR2_2534 (N9401, N9025, N8540);
not NOT1_2535 (N9402, N8541_t0);
nand NAND2_2536 (N9407, N8548_t0, N89_t0);
and AND2_2537 (N9408, N8541_t1, N8548_t1);
not NOT1_2538 (N9412, N8811_t0);
not NOT1_2539 (N9413, N8566_t0);
not NOT1_2540 (N9414, N8569_t0);
not NOT1_2541 (N9415, N8572_t0);
not NOT1_2542 (N9416, N8575_t0);
nor NOR2_2543 (N9417, N9053, N8578);
nor NOR2_2544 (N9418, N9054, N8579);
and AND3_2545 (N9419, N7387_t1, N6177_t1, N8566_t1);
and AND3_2546 (N9420, N8555_t0, N7384_t0, N8569_t1);
and AND3_2547 (N9421, N7398_t1, N7394_t1, N8572_t1);
and AND3_2548 (N9422, N8561_t0, N8558_t0, N8575_t1);
buf BUFF1_2549 (N9423, N8326_t5);
nand NAND2_2550 (N9426, N9064, N8608);
nand NAND2_2551 (N9429, N9065, N8610);
nand NAND2_2552 (N9432, N3515_t1, N9066);
nand NAND2_2553 (N9435, N4796_t1, N9072);
nand NAND2_2554 (N9442, N3628_t1, N9087);
nand NAND2_2555 (N9445, N4814_t1, N9093);
not NOT1_2556 (N9454, N8678_t0);
not NOT1_2557 (N9455, N8681_t0);
not NOT1_2558 (N9456, N8684_t0);
not NOT1_2559 (N9459, N8690_t0);
not NOT1_2560 (N9460, N8693_t0);
not NOT1_2561 (N9461, N8696_t0);
buf BUFF1_2562 (N9462, N8358_t4);
not NOT1_2563 (N9465, N8702_t0);
not NOT1_2564 (N9466, N8705_t0);
not NOT1_2565 (N9467, N8708_t0);
not NOT1_2566 (N9468, N8724_t0);
buf BUFF1_2567 (N9473, N8358_t5);
not NOT1_2568 (N9476, N8718_t0);
not NOT1_2569 (N9477, N8721_t0);
nand NAND2_2570 (N9478, N9159, N9160);
nand NAND2_2571 (N9485, N9179, N9180);
nand NAND2_2572 (N9488, N9181, N9182);
not NOT1_2573 (N9493, N8757_t0);
not NOT1_2574 (N9494, N8760_t0);
not NOT1_2575 (N9495, N8763_t0);
not NOT1_2576 (N9498, N8769_t0);
not NOT1_2577 (N9499, N8772_t0);
not NOT1_2578 (N9500, N8775_t0);
not NOT1_2579 (N9505, N8781_t0);
not NOT1_2580 (N9506, N8784_t0);
not NOT1_2581 (N9507, N8787_t0);
not NOT1_2582 (N9508, N8790_t0);
not NOT1_2583 (N9509, N8808_t0);
not NOT1_2584 (N9514, N8799_t0);
not NOT1_2585 (N9515, N8802_t0);
not NOT1_2586 (N9516, N8805_t0);
nand NAND2_2587 (N9517, N9234, N9235);
nand NAND2_2588 (N9520, N9236, N9237);
and AND2_2589 (N9526, N8943_t0, N8421_t0);
and AND2_2590 (N9531, N8943_t1, N8421_t1);
nand NAND2_2591 (N9539, N9271, N8880);
nand NAND2_2592 (N9540, N9273, N8884);
not NOT1_2593 (N9541, N9275);
and AND2_2594 (N9543, N8857_t0, N8254);
and AND2_2595 (N9551, N8871_t0, N8288);
nand NAND2_2596 (N9555, N9272, N8882);
nand NAND2_2597 (N9556, N9274, N8886);
not NOT1_2598 (N9557, N8898_t0);
and AND2_2599 (N9560, N8902_t0, N8333_t1);
not NOT1_2600 (N9561, N9099_t0);
nand NAND2_2601 (N9562, N9099_t1, N9290);
not NOT1_2602 (N9563, N9103_t0);
nand NAND2_2603 (N9564, N9103_t1, N9292);
not NOT1_2604 (N9565, N9107_t0);
nand NAND2_2605 (N9566, N9107_t1, N9294);
not NOT1_2606 (N9567, N9111_t0);
nand NAND2_2607 (N9568, N9111_t1, N9296);
nand NAND2_2608 (N9569, N4844_t1, N9298);
nand NAND2_2609 (N9570, N6207_t1, N9300);
not NOT1_2610 (N9571, N8920_t0);
not NOT1_2611 (N9575, N8927_t0);
and AND2_2612 (N9579, N8365_t1, N8927_t1);
not NOT1_2613 (N9581, N8950_t0);
not NOT1_2614 (N9582, N8956_t0);
and AND2_2615 (N9585, N8405_t2, N8956_t1);
and AND2_2616 (N9591, N8966_t0, N8430_t1);
not NOT1_2617 (N9592, N9161_t0);
nand NAND2_2618 (N9593, N9161_t1, N9352);
not NOT1_2619 (N9594, N9165_t0);
nand NAND2_2620 (N9595, N9165_t1, N9354);
not NOT1_2621 (N9596, N9169_t0);
nand NAND2_2622 (N9597, N9169_t1, N9356);
not NOT1_2623 (N9598, N9173_t0);
nand NAND2_2624 (N9599, N9173_t1, N9358);
nand NAND2_2625 (N9600, N4940_t1, N9360);
nand NAND2_2626 (N9601, N6220_t1, N9362);
and AND3_2627 (N9602, N8457_t1, N7198_t2, N9363);
and AND3_2628 (N9603, N7194_t2, N8460_t1, N9364);
and AND3_2629 (N9604, N8463_t1, N7209_t2, N9365);
and AND3_2630 (N9605, N7205_t2, N8466_t1, N9366);
not NOT1_2631 (N9608, N9001_t0);
and AND2_2632 (N9611, N8485_t1, N9001_t1);
and AND3_2633 (N9612, N8519_t1, N7318_t2, N9392);
and AND3_2634 (N9613, N7314_t2, N8522_t1, N9393);
and AND3_2635 (N9614, N7325_t1, N6131_t2, N9394);
and AND3_2636 (N9615, N6127_t2, N7328_t1, N9395);
not NOT1_2637 (N9616, N9029_t0);
not NOT1_2638 (N9617, N9035_t0);
and AND2_2639 (N9618, N8541_t2, N9035_t1);
and AND3_2640 (N9621, N7384_t1, N7387_t2, N9413);
and AND3_2641 (N9622, N6177_t2, N8555_t1, N9414);
and AND3_2642 (N9623, N8558_t1, N7398_t2, N9415);
and AND3_2643 (N9624, N7394_t2, N8561_t1, N9416);
or OR5_2644 (N9626, N4563_t1, N8352, N8353, N8354, N9285);
or OR4_2645 (N9629, N4566_t2, N8355, N8356, N9286);
or OR3_2646 (N9632, N4570_t3, N8357, N9287);
or OR2_2647 (N9635, N5960_t4, N9288);
nand NAND2_2648 (N9642, N9067, N9432);
not NOT1_2649 (N9645, N9068_t0);
nand NAND2_2650 (N9646, N9073, N9435);
not NOT1_2651 (N9649, N9074_t0);
nand NAND2_2652 (N9650, N9257, N9256);
nand NAND2_2653 (N9653, N9259, N9258);
nand NAND2_2654 (N9656, N9261, N9260);
not NOT1_2655 (N9659, N9079_t0);
nand NAND2_2656 (N9660, N9079_t1, N4809);
not NOT1_2657 (N9661, N9083_t0);
nand NAND2_2658 (N9662, N9083_t1, N6202);
nand NAND2_2659 (N9663, N9088, N9442);
not NOT1_2660 (N9666, N9089_t0);
nand NAND2_2661 (N9667, N9094, N9445);
not NOT1_2662 (N9670, N9095_t0);
or OR2_2663 (N9671, N8924_t0, N8393);
not NOT1_2664 (N9674, N9117_t0);
not NOT1_2665 (N9675, N8924_t1);
not NOT1_2666 (N9678, N9127_t0);
or OR4_2667 (N9679, N4597_t4, N8388, N8389, N9315);
or OR2_2668 (N9682, N8931_t0, N9318);
or OR5_2669 (N9685, N4593_t2, N8382, N8383, N8384, N9314);
not NOT1_2670 (N9690, N9146_t0);
nand NAND2_2671 (N9691, N9146_t1, N8717);
not NOT1_2672 (N9692, N8931_t1);
not NOT1_2673 (N9695, N9149_t0);
nand NAND2_2674 (N9698, N9401, N9400);
nand NAND2_2675 (N9702, N9368, N9367);
or OR2_2676 (N9707, N8996_t0, N8517);
not NOT1_2677 (N9710, N9183_t0);
not NOT1_2678 (N9711, N8996_t1);
not NOT1_2679 (N9714, N9193_t0);
not NOT1_2680 (N9715, N9203_t0);
nand NAND2_2681 (N9716, N9203_t1, N6235);
or OR2_2682 (N9717, N9005_t0, N8518);
not NOT1_2683 (N9720, N9206_t0);
not NOT1_2684 (N9721, N9220_t0);
nand NAND2_2685 (N9722, N9220_t1, N7573);
not NOT1_2686 (N9723, N9005_t1);
not NOT1_2687 (N9726, N9223_t0);
nand NAND2_2688 (N9727, N9418, N9417);
and AND2_2689 (N9732, N9268_t0, N8269_t0);
nand NAND2_2690 (N9733, N9581, N9326);
and AND5_2691 (N9734, N89_t1, N9408_t0, N9332_t0, N8394_t0, N8421_t2);
and AND5_2692 (N9735, N89_t2, N9408_t1, N9332_t1, N8394_t1, N8421_t3);
and AND2_2693 (N9736, N9265_t0, N8262_t0);
not NOT1_2694 (N9737, N9555);
not NOT1_2695 (N9738, N9556);
nand NAND2_2696 (N9739, N9361, N9601);
nand NAND2_2697 (N9740, N9423_t0, N1115);
not NOT1_2698 (N9741, N9423_t1);
nand NAND2_2699 (N9742, N9299, N9570);
and AND2_2700 (N9754, N8333_t2, N9280_t0);
or OR2_2701 (N9758, N8898_t1, N9560);
nand NAND2_2702 (N9762, N8660_t1, N9561);
nand NAND2_2703 (N9763, N8663_t1, N9563);
nand NAND2_2704 (N9764, N8666_t1, N9565);
nand NAND2_2705 (N9765, N8669_t1, N9567);
nand NAND2_2706 (N9766, N9297, N9569);
and AND2_2707 (N9767, N9280_t1, N367_t6);
nand NAND2_2708 (N9768, N9557, N9276);
not NOT1_2709 (N9769, N9307_t0);
nand NAND2_2710 (N9773, N9307_t1, N367_t7);
nand NAND2_2711 (N9774, N9571, N9301);
and AND2_2712 (N9775, N8365_t2, N9307_t2);
or OR2_2713 (N9779, N8920_t1, N9579);
not NOT1_2714 (N9784, N9478_t0);
nand NAND2_2715 (N9785, N9616, N9402);
or OR2_2716 (N9786, N8950_t1, N9585);
and AND4_2717 (N9790, N89_t3, N9408_t2, N9332_t2, N8394_t2);
or OR2_2718 (N9791, N8963, N9591);
nand NAND2_2719 (N9795, N8735_t1, N9592);
nand NAND2_2720 (N9796, N8738_t1, N9594);
nand NAND2_2721 (N9797, N8741_t1, N9596);
nand NAND2_2722 (N9798, N8744_t1, N9598);
nand NAND2_2723 (N9799, N9359, N9600);
nor NOR2_2724 (N9800, N9602, N9369);
nor NOR2_2725 (N9801, N9603, N9370);
nor NOR2_2726 (N9802, N9604, N9371);
nor NOR2_2727 (N9803, N9605, N9372);
not NOT1_2728 (N9805, N9485_t0);
not NOT1_2729 (N9806, N9488_t0);
or OR2_2730 (N9809, N8995, N9611);
nor NOR2_2731 (N9813, N9612, N9396);
nor NOR2_2732 (N9814, N9613, N9397);
nor NOR2_2733 (N9815, N9614, N9398);
nor NOR2_2734 (N9816, N9615, N9399);
and AND2_2735 (N9817, N9617, N9407);
or OR2_2736 (N9820, N9029_t1, N9618);
not NOT1_2737 (N9825, N9517_t0);
not NOT1_2738 (N9826, N9520_t0);
nor NOR2_2739 (N9827, N9621, N9419);
nor NOR2_2740 (N9828, N9622, N9420);
nor NOR2_2741 (N9829, N9623, N9421);
nor NOR2_2742 (N9830, N9624, N9422);
not NOT1_2743 (N9835, N9426_t0);
nand NAND2_2744 (N9836, N9426_t1, N4789);
not NOT1_2745 (N9837, N9429_t0);
nand NAND2_2746 (N9838, N9429_t1, N4794);
nand NAND2_2747 (N9846, N3625_t1, N9659);
nand NAND2_2748 (N9847, N4810_t1, N9661);
not NOT1_2749 (N9862, N9462_t0);
nand NAND2_2750 (N9863, N7553_t1, N9690);
not NOT1_2751 (N9866, N9473_t0);
nand NAND2_2752 (N9873, N5030_t1, N9715);
nand NAND2_2753 (N9876, N6236_t1, N9721);
nand NAND2_2754 (N9890, N9795, N9593);
nand NAND2_2755 (N9891, N9797, N9597);
not NOT1_2756 (N9892, N9799);
nand NAND2_2757 (N9893, N871_t1, N9741);
nand NAND2_2758 (N9894, N9762, N9562);
nand NAND2_2759 (N9895, N9764, N9566);
not NOT1_2760 (N9896, N9766);
not NOT1_2761 (N9897, N9626_t0);
nand NAND2_2762 (N9898, N9626_t1, N9249);
not NOT1_2763 (N9899, N9629_t0);
nand NAND2_2764 (N9900, N9629_t1, N9250);
not NOT1_2765 (N9901, N9632_t0);
nand NAND2_2766 (N9902, N9632_t1, N9251);
not NOT1_2767 (N9903, N9635_t0);
nand NAND2_2768 (N9904, N9635_t1, N9252);
not NOT1_2769 (N9905, N9543_t0);
not NOT1_2770 (N9906, N9650_t0);
nand NAND2_2771 (N9907, N9650_t1, N5769);
not NOT1_2772 (N9908, N9653_t0);
nand NAND2_2773 (N9909, N9653_t1, N5770);
not NOT1_2774 (N9910, N9656_t0);
nand NAND2_2775 (N9911, N9656_t1, N9262);
not NOT1_2776 (N9917, N9551_t0);
nand NAND2_2777 (N9923, N9763, N9564);
nand NAND2_2778 (N9924, N9765, N9568);
or OR2_2779 (N9925, N8902_t1, N9767);
and AND2_2780 (N9932, N9575_t0, N9773);
and AND2_2781 (N9935, N9575_t1, N9769);
not NOT1_2782 (N9938, N9698_t0);
nand NAND2_2783 (N9939, N9698_t1, N9323);
nand NAND2_2784 (N9945, N9796, N9595);
nand NAND2_2785 (N9946, N9798, N9599);
not NOT1_2786 (N9947, N9702_t0);
nand NAND2_2787 (N9948, N9702_t1, N6102);
and AND2_2788 (N9949, N9608_t0, N9375);
not NOT1_2789 (N9953, N9727_t0);
nand NAND2_2790 (N9954, N9727_t1, N9412);
nand NAND2_2791 (N9955, N3502_t1, N9835);
nand NAND2_2792 (N9956, N3510_t1, N9837);
not NOT1_2793 (N9957, N9642_t0);
nand NAND2_2794 (N9958, N9642_t1, N9645);
not NOT1_2795 (N9959, N9646_t0);
nand NAND2_2796 (N9960, N9646_t1, N9649);
nand NAND2_2797 (N9961, N9660, N9846);
nand NAND2_2798 (N9964, N9662, N9847);
not NOT1_2799 (N9967, N9663_t0);
nand NAND2_2800 (N9968, N9663_t1, N9666);
not NOT1_2801 (N9969, N9667_t0);
nand NAND2_2802 (N9970, N9667_t1, N9670);
not NOT1_2803 (N9971, N9671_t0);
nand NAND2_2804 (N9972, N9671_t1, N6213);
not NOT1_2805 (N9973, N9675_t0);
nand NAND2_2806 (N9974, N9675_t1, N7551);
not NOT1_2807 (N9975, N9679_t0);
nand NAND2_2808 (N9976, N9679_t1, N7552);
not NOT1_2809 (N9977, N9682_t0);
not NOT1_2810 (N9978, N9685_t0);
nand NAND2_2811 (N9979, N9691, N9863);
not NOT1_2812 (N9982, N9692_t0);
nand NAND2_2813 (N9983, N9814, N9813);
nand NAND2_2814 (N9986, N9816, N9815);
nand NAND2_2815 (N9989, N9801, N9800);
nand NAND2_2816 (N9992, N9803, N9802);
not NOT1_2817 (N9995, N9707_t0);
nand NAND2_2818 (N9996, N9707_t1, N6231);
not NOT1_2819 (N9997, N9711_t0);
nand NAND2_2820 (N9998, N9711_t1, N7572);
nand NAND2_2821 (N9999, N9716, N9873);
not NOT1_2822 (N10002, N9717_t0);
nand NAND2_2823 (N10003, N9722, N9876);
not NOT1_2824 (N10006, N9723_t0);
nand NAND2_2825 (N10007, N9830, N9829);
nand NAND2_2826 (N10010, N9828, N9827);
and AND3_2827 (N10013, N9791_t0, N8307_t0, N8269_t1);
and AND4_2828 (N10014, N9758_t0, N9344_t0, N8307_t1, N8269_t2);
and AND5_2829 (N10015, N367_t8, N9754_t0, N9344_t1, N8307_t2, N8269_t3);
and AND3_2830 (N10016, N9786_t0, N8394_t3, N8421_t4);
and AND4_2831 (N10017, N9820_t0, N9332_t3, N8394_t4, N8421_t5);
and AND3_2832 (N10018, N9786_t1, N8394_t5, N8421_t6);
and AND4_2833 (N10019, N9820_t1, N9332_t4, N8394_t6, N8421_t7);
and AND3_2834 (N10020, N9809_t0, N8298_t0, N8262_t1);
and AND4_2835 (N10021, N9779_t0, N9385_t0, N8298_t1, N8262_t2);
and AND5_2836 (N10022, N367_t9, N9775_t0, N9385_t1, N8298_t2, N8262_t3);
not NOT1_2837 (N10023, N9945);
not NOT1_2838 (N10024, N9946);
nand NAND2_2839 (N10025, N9740, N9893);
not NOT1_2840 (N10026, N9923);
not NOT1_2841 (N10028, N9924);
nand NAND2_2842 (N10032, N8595_t1, N9897);
nand NAND2_2843 (N10033, N8598_t1, N9899);
nand NAND2_2844 (N10034, N8601_t1, N9901);
nand NAND2_2845 (N10035, N8604_t1, N9903);
nand NAND2_2846 (N10036, N4803_t1, N9906);
nand NAND2_2847 (N10037, N4806_t1, N9908);
nand NAND2_2848 (N10038, N8627_t1, N9910);
and AND2_2849 (N10039, N9809_t1, N8298_t3);
and AND3_2850 (N10040, N9779_t1, N9385_t2, N8298_t4);
and AND4_2851 (N10041, N367_t10, N9775_t1, N9385_t3, N8298_t5);
and AND2_2852 (N10042, N9779_t2, N9385_t4);
and AND3_2853 (N10043, N367_t11, N9775_t2, N9385_t5);
nand NAND2_2854 (N10050, N8727_t1, N9938);
not NOT1_2855 (N10053, N9817_t0);
and AND2_2856 (N10054, N9817_t1, N9029_t2);
and AND2_2857 (N10055, N9786_t2, N8394_t7);
and AND3_2858 (N10056, N9820_t2, N9332_t5, N8394_t8);
and AND2_2859 (N10057, N9791_t1, N8307_t3);
and AND3_2860 (N10058, N9758_t1, N9344_t2, N8307_t4);
and AND4_2861 (N10059, N367_t12, N9754_t1, N9344_t3, N8307_t5);
and AND2_2862 (N10060, N9758_t2, N9344_t4);
and AND3_2863 (N10061, N367_t13, N9754_t2, N9344_t5);
nand NAND2_2864 (N10062, N4997_t1, N9947);
nand NAND2_2865 (N10067, N8811_t1, N9953);
nand NAND2_2866 (N10070, N9955, N9836);
nand NAND2_2867 (N10073, N9956, N9838);
nand NAND2_2868 (N10076, N9068_t1, N9957);
nand NAND2_2869 (N10077, N9074_t1, N9959);
nand NAND2_2870 (N10082, N9089_t1, N9967);
nand NAND2_2871 (N10083, N9095_t1, N9969);
nand NAND2_2872 (N10084, N4871_t1, N9971);
nand NAND2_2873 (N10085, N6214_t1, N9973);
nand NAND2_2874 (N10086, N6217_t1, N9975);
nand NAND2_2875 (N10093, N5027_t1, N9995);
nand NAND2_2876 (N10094, N6232_t1, N9997);
or OR5_2877 (N10101, N9238, N9732, N10013, N10014, N10015);
or OR5_2878 (N10102, N9339_t0, N9526, N10016, N10017, N9734);
or OR5_2879 (N10103, N9339_t1, N9531, N10018, N10019, N9735);
or OR5_2880 (N10104, N9242, N9736, N10020, N10021, N10022);
and AND2_2881 (N10105, N9925_t0, N9894);
and AND2_2882 (N10106, N9925_t1, N9895);
and AND2_2883 (N10107, N9925_t2, N9896);
and AND2_2884 (N10108, N9925_t3, N8253);
nand NAND2_2885 (N10109, N10032, N9898);
nand NAND2_2886 (N10110, N10033, N9900);
nand NAND2_2887 (N10111, N10034, N9902);
nand NAND2_2888 (N10112, N10035, N9904);
nand NAND2_2889 (N10113, N10036, N9907);
nand NAND2_2890 (N10114, N10037, N9909);
nand NAND2_2891 (N10115, N10038, N9911);
or OR4_2892 (N10116, N9265_t1, N10039, N10040, N10041);
or OR3_2893 (N10119, N9809_t2, N10042, N10043);
not NOT1_2894 (N10124, N9925_t4);
and AND2_2895 (N10130, N9768, N9925_t5);
not NOT1_2896 (N10131, N9932_t0);
not NOT1_2897 (N10132, N9935_t0);
and AND2_2898 (N10133, N9932_t1, N8920_t2);
nand NAND2_2899 (N10134, N10050, N9939);
not NOT1_2900 (N10135, N9983_t0);
nand NAND2_2901 (N10136, N9983_t1, N9324);
not NOT1_2902 (N10137, N9986_t0);
nand NAND2_2903 (N10138, N9986_t1, N9784);
and AND2_2904 (N10139, N9785, N10053);
or OR4_2905 (N10140, N8943_t2, N10055, N10056, N9790);
or OR4_2906 (N10141, N9268_t1, N10057, N10058, N10059);
or OR3_2907 (N10148, N9791_t2, N10060, N10061);
nand NAND2_2908 (N10155, N10062, N9948);
not NOT1_2909 (N10156, N9989_t0);
nand NAND2_2910 (N10157, N9989_t1, N9805);
not NOT1_2911 (N10158, N9992_t0);
nand NAND2_2912 (N10159, N9992_t1, N9806);
not NOT1_2913 (N10160, N9949_t0);
nand NAND2_2914 (N10161, N10067, N9954);
not NOT1_2915 (N10162, N10007_t0);
nand NAND2_2916 (N10163, N10007_t1, N9825);
not NOT1_2917 (N10164, N10010_t0);
nand NAND2_2918 (N10165, N10010_t1, N9826);
nand NAND2_2919 (N10170, N10076, N9958);
nand NAND2_2920 (N10173, N10077, N9960);
not NOT1_2921 (N10176, N9961_t0);
nand NAND2_2922 (N10177, N9961_t1, N9082);
not NOT1_2923 (N10178, N9964_t0);
nand NAND2_2924 (N10179, N9964_t1, N9086);
nand NAND2_2925 (N10180, N10082, N9968);
nand NAND2_2926 (N10183, N10083, N9970);
nand NAND2_2927 (N10186, N9972, N10084);
nand NAND2_2928 (N10189, N9974, N10085);
nand NAND2_2929 (N10192, N9976, N10086);
not NOT1_2930 (N10195, N9979_t0);
nand NAND2_2931 (N10196, N9979_t1, N9982);
nand NAND2_2932 (N10197, N9996, N10093);
nand NAND2_2933 (N10200, N9998, N10094);
not NOT1_2934 (N10203, N9999_t0);
nand NAND2_2935 (N10204, N9999_t1, N10002);
not NOT1_2936 (N10205, N10003_t0);
nand NAND2_2937 (N10206, N10003_t1, N10006);
nand NAND2_2938 (N10212, N10070_t0, N4308);
nand NAND2_2939 (N10213, N10073_t0, N4313);
and AND2_2940 (N10230, N9774, N10131);
nand NAND2_2941 (N10231, N8730_t1, N10135);
nand NAND2_2942 (N10232, N9478_t1, N10137);
or OR2_2943 (N10233, N10139, N10054);
nand NAND2_2944 (N10234, N7100_t1, N10140);
nand NAND2_2945 (N10237, N9485_t1, N10156);
nand NAND2_2946 (N10238, N9488_t1, N10158);
nand NAND2_2947 (N10239, N9517_t1, N10162);
nand NAND2_2948 (N10240, N9520_t1, N10164);
not NOT1_2949 (N10241, N10070_t1);
not NOT1_2950 (N10242, N10073_t1);
nand NAND2_2951 (N10247, N8146_t1, N10176);
nand NAND2_2952 (N10248, N8156_t1, N10178);
nand NAND2_2953 (N10259, N9692_t1, N10195);
nand NAND2_2954 (N10264, N9717_t1, N10203);
nand NAND2_2955 (N10265, N9723_t1, N10205);
and AND2_2956 (N10266, N10026, N10124_t0);
and AND2_2957 (N10267, N10028, N10124_t1);
and AND2_2958 (N10268, N9742, N10124_t2);
and AND2_2959 (N10269, N6923_t4, N10124_t3);
nand NAND2_2960 (N10270, N6762_t2, N10116_t0);
nand NAND2_2961 (N10271, N3061_t1, N10241);
nand NAND2_2962 (N10272, N3064_t1, N10242);
buf BUFF1_2963 (N10273, N10116_t1);
and AND5_2964 (N10278, N10141_t0, N5728_t2, N5707_t8, N5718_t6, N5697_t8);
and AND4_2965 (N10279, N10141_t1, N5728_t3, N5707_t9, N5718_t7);
and AND3_2966 (N10280, N10141_t2, N5728_t4, N5718_t8);
and AND2_2967 (N10281, N10141_t3, N5728_t5);
and AND2_2968 (N10282, N6784_t1, N10141_t4);
not NOT1_2969 (N10283, N10119_t0);
and AND5_2970 (N10287, N10148_t0, N5936_t2, N5915_t8, N5926_t6, N5905_t8);
and AND4_2971 (N10288, N10148_t1, N5936_t3, N5915_t9, N5926_t7);
and AND3_2972 (N10289, N10148_t2, N5936_t4, N5926_t8);
and AND2_2973 (N10290, N10148_t3, N5936_t5);
and AND2_2974 (N10291, N6881_t1, N10148_t4);
and AND2_2975 (N10292, N8898_t2, N10124_t4);
nand NAND2_2976 (N10293, N10231, N10136);
nand NAND2_2977 (N10294, N10232, N10138);
nand NAND2_2978 (N10295, N8412_t1, N10233);
and AND2_2979 (N10296, N8959, N10234);
nand NAND2_2980 (N10299, N10237, N10157);
nand NAND2_2981 (N10300, N10238, N10159);
or OR2_2982 (N10301, N10230, N10133);
nand NAND2_2983 (N10306, N10239, N10163);
nand NAND2_2984 (N10307, N10240, N10165);
buf BUFF1_2985 (N10308, N10148_t5);
buf BUFF1_2986 (N10311, N10141_t5);
not NOT1_2987 (N10314, N10170_t0);
nand NAND2_2988 (N10315, N10170_t1, N9071);
not NOT1_2989 (N10316, N10173_t0);
nand NAND2_2990 (N10317, N10173_t1, N9077);
nand NAND2_2991 (N10318, N10247, N10177);
nand NAND2_2992 (N10321, N10248, N10179);
not NOT1_2993 (N10324, N10180_t0);
nand NAND2_2994 (N10325, N10180_t1, N9092);
not NOT1_2995 (N10326, N10183_t0);
nand NAND2_2996 (N10327, N10183_t1, N9098);
not NOT1_2997 (N10328, N10186_t0);
nand NAND2_2998 (N10329, N10186_t1, N9674);
not NOT1_2999 (N10330, N10189_t0);
nand NAND2_3000 (N10331, N10189_t1, N9678);
not NOT1_3001 (N10332, N10192_t0);
nand NAND2_3002 (N10333, N10192_t1, N9977);
nand NAND2_3003 (N10334, N10259, N10196);
not NOT1_3004 (N10337, N10197_t0);
nand NAND2_3005 (N10338, N10197_t1, N9710);
not NOT1_3006 (N10339, N10200_t0);
nand NAND2_3007 (N10340, N10200_t1, N9714);
nand NAND2_3008 (N10341, N10264, N10204);
nand NAND2_3009 (N10344, N10265, N10206);
or OR2_3010 (N10350, N10266, N10105);
or OR2_3011 (N10351, N10267, N10106);
or OR2_3012 (N10352, N10268, N10107);
or OR2_3013 (N10353, N10269, N10108);
and AND2_3014 (N10354, N8857_t1, N10270);
nand NAND2_3015 (N10357, N10271, N10212);
nand NAND2_3016 (N10360, N10272, N10213);
or OR2_3017 (N10367, N7620_t1, N10282);
or OR2_3018 (N10375, N7671_t1, N10291);
or OR2_3019 (N10381, N10292, N10130);
and AND4_3020 (N10388, N10114, N10134, N10293, N10294);
and AND2_3021 (N10391, N9582, N10295);
and AND4_3022 (N10399, N10113, N10115, N10299, N10300);
and AND4_3023 (N10402, N10155, N10161, N10306, N10307);
or OR5_3024 (N10406, N3229_t1, N6888, N6889, N6890, N10287);
or OR4_3025 (N10409, N3232_t2, N6891, N6892, N10288);
or OR3_3026 (N10412, N3236_t3, N6893, N10289);
or OR2_3027 (N10415, N3241_t4, N10290);
or OR5_3028 (N10419, N3137_t1, N6791, N6792, N6793, N10278);
or OR4_3029 (N10422, N3140_t2, N6794, N6795, N10279);
or OR3_3030 (N10425, N3144_t3, N6796, N10280);
or OR2_3031 (N10428, N3149_t4, N10281);
nand NAND2_3032 (N10431, N8117_t1, N10314);
nand NAND2_3033 (N10432, N8134_t1, N10316);
nand NAND2_3034 (N10437, N8169_t1, N10324);
nand NAND2_3035 (N10438, N8186_t1, N10326);
nand NAND2_3036 (N10439, N9117_t1, N10328);
nand NAND2_3037 (N10440, N9127_t1, N10330);
nand NAND2_3038 (N10441, N9682_t1, N10332);
nand NAND2_3039 (N10444, N9183_t1, N10337);
nand NAND2_3040 (N10445, N9193_t1, N10339);
not NOT1_3041 (N10450, N10296_t0);
and AND2_3042 (N10451, N10296_t1, N4193_t2);
not NOT1_3043 (N10455, N10308_t0);
nand NAND2_3044 (N10456, N10308_t1, N8242);
not NOT1_3045 (N10465, N10311_t0);
nand NAND2_3046 (N10466, N10311_t1, N8247);
not NOT1_3047 (N10479, N10273_t0);
not NOT1_3048 (N10497, N10301_t0);
nand NAND2_3049 (N10509, N10431, N10315);
nand NAND2_3050 (N10512, N10432, N10317);
not NOT1_3051 (N10515, N10318_t0);
nand NAND2_3052 (N10516, N10318_t1, N8632);
not NOT1_3053 (N10517, N10321_t0);
nand NAND2_3054 (N10518, N10321_t1, N8637);
nand NAND2_3055 (N10519, N10437, N10325);
nand NAND2_3056 (N10522, N10438, N10327);
nand NAND2_3057 (N10525, N10439, N10329);
nand NAND2_3058 (N10528, N10440, N10331);
nand NAND2_3059 (N10531, N10441, N10333);
not NOT1_3060 (N10534, N10334_t0);
nand NAND2_3061 (N10535, N10334_t1, N9695);
nand NAND2_3062 (N10536, N10444, N10338);
nand NAND2_3063 (N10539, N10445, N10340);
not NOT1_3064 (N10542, N10341_t0);
nand NAND2_3065 (N10543, N10341_t1, N9720);
not NOT1_3066 (N10544, N10344_t0);
nand NAND2_3067 (N10545, N10344_t1, N9726);
and AND2_3068 (N10546, N5631, N10450);
not NOT1_3069 (N10547, N10391_t0);
and AND2_3070 (N10548, N10391_t1, N8950_t2);
and AND2_3071 (N10549, N5165, N10367_t0);
not NOT1_3072 (N10550, N10354_t0);
and AND2_3073 (N10551, N10354_t1, N3126_t2);
nand NAND2_3074 (N10552, N7411_t1, N10455);
and AND2_3075 (N10553, N10375_t0, N9539);
and AND2_3076 (N10554, N10375_t1, N9540);
and AND2_3077 (N10555, N10375_t2, N9541);
and AND2_3078 (N10556, N10375_t3, N6761);
not NOT1_3079 (N10557, N10406_t0);
nand NAND2_3080 (N10558, N10406_t1, N8243);
not NOT1_3081 (N10559, N10409_t0);
nand NAND2_3082 (N10560, N10409_t1, N8244);
not NOT1_3083 (N10561, N10412_t0);
nand NAND2_3084 (N10562, N10412_t1, N8245);
not NOT1_3085 (N10563, N10415_t0);
nand NAND2_3086 (N10564, N10415_t1, N8246);
nand NAND2_3087 (N10565, N7426_t1, N10465);
not NOT1_3088 (N10566, N10419_t0);
nand NAND2_3089 (N10567, N10419_t1, N8248);
not NOT1_3090 (N10568, N10422_t0);
nand NAND2_3091 (N10569, N10422_t1, N8249);
not NOT1_3092 (N10570, N10425_t0);
nand NAND2_3093 (N10571, N10425_t1, N8250);
not NOT1_3094 (N10572, N10428_t0);
nand NAND2_3095 (N10573, N10428_t1, N8251);
not NOT1_3096 (N10574, N10399_t0);
not NOT1_3097 (N10575, N10402_t0);
not NOT1_3098 (N10576, N10388_t0);
and AND3_3099 (N10577, N10399_t1, N10402_t1, N10388_t1);
and AND3_3100 (N10581, N10360_t0, N9543_t1, N10273_t1);
and AND3_3101 (N10582, N10357_t0, N9905, N10273_t2);
not NOT1_3102 (N10583, N10367_t1);
and AND2_3103 (N10587, N10367_t2, N5735);
and AND2_3104 (N10588, N10367_t3, N3135);
not NOT1_3105 (N10589, N10375_t4);
and AND5_3106 (N10594, N10381_t0, N7180_t2, N7159_t8, N7170_t6, N7149_t8);
and AND4_3107 (N10595, N10381_t1, N7180_t3, N7159_t9, N7170_t7);
and AND3_3108 (N10596, N10381_t2, N7180_t4, N7170_t8);
and AND2_3109 (N10597, N10381_t3, N7180_t5);
and AND2_3110 (N10598, N8444_t1, N10381_t4);
buf BUFF1_3111 (N10602, N10381_t5);
nand NAND2_3112 (N10609, N7479_t1, N10515);
nand NAND2_3113 (N10610, N7491_t1, N10517);
nand NAND2_3114 (N10621, N9149_t1, N10534);
nand NAND2_3115 (N10626, N9206_t1, N10542);
nand NAND2_3116 (N10627, N9223_t1, N10544);
or OR2_3117 (N10628, N10546, N10451);
and AND2_3118 (N10629, N9733, N10547);
and AND2_3119 (N10631, N5166, N10550);
nand NAND2_3120 (N10632, N10552, N10456);
nand NAND2_3121 (N10637, N7414_t1, N10557);
nand NAND2_3122 (N10638, N7417_t1, N10559);
nand NAND2_3123 (N10639, N7420_t1, N10561);
nand NAND2_3124 (N10640, N7423_t1, N10563);
nand NAND2_3125 (N10641, N10565, N10466);
nand NAND2_3126 (N10642, N7429_t1, N10566);
nand NAND2_3127 (N10643, N7432_t1, N10568);
nand NAND2_3128 (N10644, N7435_t1, N10570);
nand NAND2_3129 (N10645, N7438_t1, N10572);
and AND3_3130 (N10647, N886, N887, N10577);
and AND3_3131 (N10648, N10360_t1, N8857_t2, N10479_t0);
and AND3_3132 (N10649, N10357_t1, N7609_t2, N10479_t1);
or OR2_3133 (N10652, N8966_t1, N10598);
or OR5_3134 (N10659, N4675_t1, N8451, N8452, N8453, N10594);
or OR4_3135 (N10662, N4678_t2, N8454, N8455, N10595);
or OR3_3136 (N10665, N4682_t3, N8456, N10596);
or OR2_3137 (N10668, N4687_t4, N10597);
not NOT1_3138 (N10671, N10509_t0);
nand NAND2_3139 (N10672, N10509_t1, N8615);
not NOT1_3140 (N10673, N10512_t0);
nand NAND2_3141 (N10674, N10512_t1, N8624);
nand NAND2_3142 (N10675, N10609, N10516);
nand NAND2_3143 (N10678, N10610, N10518);
not NOT1_3144 (N10681, N10519_t0);
nand NAND2_3145 (N10682, N10519_t1, N8644);
not NOT1_3146 (N10683, N10522_t0);
nand NAND2_3147 (N10684, N10522_t1, N8653);
not NOT1_3148 (N10685, N10525_t0);
nand NAND2_3149 (N10686, N10525_t1, N9454);
not NOT1_3150 (N10687, N10528_t0);
nand NAND2_3151 (N10688, N10528_t1, N9459);
not NOT1_3152 (N10689, N10531_t0);
nand NAND2_3153 (N10690, N10531_t1, N9978);
nand NAND2_3154 (N10691, N10621, N10535);
not NOT1_3155 (N10694, N10536_t0);
nand NAND2_3156 (N10695, N10536_t1, N9493);
not NOT1_3157 (N10696, N10539_t0);
nand NAND2_3158 (N10697, N10539_t1, N9498);
nand NAND2_3159 (N10698, N10626, N10543);
nand NAND2_3160 (N10701, N10627, N10545);
or OR2_3161 (N10704, N10629, N10548);
and AND2_3162 (N10705, N3159_t2, N10583_t0);
or OR2_3163 (N10706, N10631, N10551);
and AND2_3164 (N10707, N9737, N10589_t0);
and AND2_3165 (N10708, N9738, N10589_t1);
and AND2_3166 (N10709, N9243, N10589_t2);
and AND2_3167 (N10710, N5892_t4, N10589_t3);
nand NAND2_3168 (N10711, N10637, N10558);
nand NAND2_3169 (N10712, N10638, N10560);
nand NAND2_3170 (N10713, N10639, N10562);
nand NAND2_3171 (N10714, N10640, N10564);
nand NAND2_3172 (N10715, N10642, N10567);
nand NAND2_3173 (N10716, N10643, N10569);
nand NAND2_3174 (N10717, N10644, N10571);
nand NAND2_3175 (N10718, N10645, N10573);
not NOT1_3176 (N10719, N10602_t0);
nand NAND2_3177 (N10720, N10602_t1, N9244);
not NOT1_3178 (N10729, N10647);
and AND2_3179 (N10730, N5178, N10583_t1);
and AND2_3180 (N10731, N2533_t2, N10583_t2);
nand NAND2_3181 (N10737, N7447_t1, N10671);
nand NAND2_3182 (N10738, N7465_t1, N10673);
or OR4_3183 (N10739, N10648, N10649, N10581, N10582);
nand NAND2_3184 (N10746, N7503_t1, N10681);
nand NAND2_3185 (N10747, N7521_t1, N10683);
nand NAND2_3186 (N10748, N8678_t1, N10685);
nand NAND2_3187 (N10749, N8690_t1, N10687);
nand NAND2_3188 (N10750, N9685_t1, N10689);
nand NAND2_3189 (N10753, N8757_t1, N10694);
nand NAND2_3190 (N10754, N8769_t1, N10696);
or OR2_3191 (N10759, N10705, N10549);
or OR2_3192 (N10760, N10707, N10553);
or OR2_3193 (N10761, N10708, N10554);
or OR2_3194 (N10762, N10709, N10555);
or OR2_3195 (N10763, N10710, N10556);
nand NAND2_3196 (N10764, N8580_t1, N10719);
and AND2_3197 (N10765, N10652_t0, N9890);
and AND2_3198 (N10766, N10652_t1, N9891);
and AND2_3199 (N10767, N10652_t2, N9892);
and AND2_3200 (N10768, N10652_t3, N8252);
not NOT1_3201 (N10769, N10659_t0);
nand NAND2_3202 (N10770, N10659_t1, N9245);
not NOT1_3203 (N10771, N10662_t0);
nand NAND2_3204 (N10772, N10662_t1, N9246);
not NOT1_3205 (N10773, N10665_t0);
nand NAND2_3206 (N10774, N10665_t1, N9247);
not NOT1_3207 (N10775, N10668_t0);
nand NAND2_3208 (N10776, N10668_t1, N9248);
or OR2_3209 (N10778, N10730, N10587);
or OR2_3210 (N10781, N10731, N10588);
not NOT1_3211 (N10784, N10652_t4);
nand NAND2_3212 (N10789, N10737, N10672);
nand NAND2_3213 (N10792, N10738, N10674);
not NOT1_3214 (N10796, N10675_t0);
nand NAND2_3215 (N10797, N10675_t1, N8633);
not NOT1_3216 (N10798, N10678_t0);
nand NAND2_3217 (N10799, N10678_t1, N8638);
nand NAND2_3218 (N10800, N10746, N10682);
nand NAND2_3219 (N10803, N10747, N10684);
nand NAND2_3220 (N10806, N10748, N10686);
nand NAND2_3221 (N10809, N10749, N10688);
nand NAND2_3222 (N10812, N10750, N10690);
not NOT1_3223 (N10815, N10691_t0);
nand NAND2_3224 (N10816, N10691_t1, N9866);
nand NAND2_3225 (N10817, N10753, N10695);
nand NAND2_3226 (N10820, N10754, N10697);
not NOT1_3227 (N10823, N10698_t0);
nand NAND2_3228 (N10824, N10698_t1, N9505);
not NOT1_3229 (N10825, N10701_t0);
nand NAND2_3230 (N10826, N10701_t1, N9514);
nand NAND2_3231 (N10827, N10764, N10720);
nand NAND2_3232 (N10832, N8583_t1, N10769);
nand NAND2_3233 (N10833, N8586_t1, N10771);
nand NAND2_3234 (N10834, N8589_t1, N10773);
nand NAND2_3235 (N10835, N8592_t1, N10775);
not NOT1_3236 (N10836, N10739_t0);
buf BUFF1_3237 (N10837, N10778_t0);
buf BUFF1_3238 (N10838, N10778_t1);
buf BUFF1_3239 (N10839, N10781_t0);
buf BUFF1_3240 (N10840, N10781_t1);
nand NAND2_3241 (N10845, N7482_t1, N10796);
nand NAND2_3242 (N10846, N7494_t1, N10798);
nand NAND2_3243 (N10857, N9473_t1, N10815);
nand NAND2_3244 (N10862, N8781_t1, N10823);
nand NAND2_3245 (N10863, N8799_t1, N10825);
and AND2_3246 (N10864, N10023, N10784_t0);
and AND2_3247 (N10865, N10024, N10784_t1);
and AND2_3248 (N10866, N9739, N10784_t2);
and AND2_3249 (N10867, N7136_t4, N10784_t3);
nand NAND2_3250 (N10868, N10832, N10770);
nand NAND2_3251 (N10869, N10833, N10772);
nand NAND2_3252 (N10870, N10834, N10774);
nand NAND2_3253 (N10871, N10835, N10776);
not NOT1_3254 (N10872, N10789_t0);
nand NAND2_3255 (N10873, N10789_t1, N8616);
not NOT1_3256 (N10874, N10792_t0);
nand NAND2_3257 (N10875, N10792_t1, N8625);
nand NAND2_3258 (N10876, N10845, N10797);
nand NAND2_3259 (N10879, N10846, N10799);
not NOT1_3260 (N10882, N10800_t0);
nand NAND2_3261 (N10883, N10800_t1, N8645);
not NOT1_3262 (N10884, N10803_t0);
nand NAND2_3263 (N10885, N10803_t1, N8654);
not NOT1_3264 (N10886, N10806_t0);
nand NAND2_3265 (N10887, N10806_t1, N9455);
not NOT1_3266 (N10888, N10809_t0);
nand NAND2_3267 (N10889, N10809_t1, N9460);
not NOT1_3268 (N10890, N10812_t0);
nand NAND2_3269 (N10891, N10812_t1, N9862);
nand NAND2_3270 (N10892, N10857, N10816);
not NOT1_3271 (N10895, N10817_t0);
nand NAND2_3272 (N10896, N10817_t1, N9494);
not NOT1_3273 (N10897, N10820_t0);
nand NAND2_3274 (N10898, N10820_t1, N9499);
nand NAND2_3275 (N10899, N10862, N10824);
nand NAND2_3276 (N10902, N10863, N10826);
or OR2_3277 (N10905, N10864, N10765);
or OR2_3278 (N10906, N10865, N10766);
or OR2_3279 (N10907, N10866, N10767);
or OR2_3280 (N10908, N10867, N10768);
nand NAND2_3281 (N10909, N7450_t1, N10872);
nand NAND2_3282 (N10910, N7468_t1, N10874);
nand NAND2_3283 (N10915, N7506_t1, N10882);
nand NAND2_3284 (N10916, N7524_t1, N10884);
nand NAND2_3285 (N10917, N8681_t1, N10886);
nand NAND2_3286 (N10918, N8693_t1, N10888);
nand NAND2_3287 (N10919, N9462_t1, N10890);
nand NAND2_3288 (N10922, N8760_t1, N10895);
nand NAND2_3289 (N10923, N8772_t1, N10897);
nand NAND2_3290 (N10928, N10909, N10873);
nand NAND2_3291 (N10931, N10910, N10875);
not NOT1_3292 (N10934, N10876_t0);
nand NAND2_3293 (N10935, N10876_t1, N8634);
not NOT1_3294 (N10936, N10879_t0);
nand NAND2_3295 (N10937, N10879_t1, N8639);
nand NAND2_3296 (N10938, N10915, N10883);
nand NAND2_3297 (N10941, N10916, N10885);
nand NAND2_3298 (N10944, N10917, N10887);
nand NAND2_3299 (N10947, N10918, N10889);
nand NAND2_3300 (N10950, N10919, N10891);
not NOT1_3301 (N10953, N10892_t0);
nand NAND2_3302 (N10954, N10892_t1, N9476);
nand NAND2_3303 (N10955, N10922, N10896);
nand NAND2_3304 (N10958, N10923, N10898);
not NOT1_3305 (N10961, N10899_t0);
nand NAND2_3306 (N10962, N10899_t1, N9506);
not NOT1_3307 (N10963, N10902_t0);
nand NAND2_3308 (N10964, N10902_t1, N9515);
nand NAND2_3309 (N10969, N7485_t1, N10934);
nand NAND2_3310 (N10970, N7497_t1, N10936);
nand NAND2_3311 (N10981, N8718_t1, N10953);
nand NAND2_3312 (N10986, N8784_t1, N10961);
nand NAND2_3313 (N10987, N8802_t1, N10963);
not NOT1_3314 (N10988, N10928_t0);
nand NAND2_3315 (N10989, N10928_t1, N8617);
not NOT1_3316 (N10990, N10931_t0);
nand NAND2_3317 (N10991, N10931_t1, N8626);
nand NAND2_3318 (N10992, N10969, N10935);
nand NAND2_3319 (N10995, N10970, N10937);
not NOT1_3320 (N10998, N10938_t0);
nand NAND2_3321 (N10999, N10938_t1, N8646);
not NOT1_3322 (N11000, N10941_t0);
nand NAND2_3323 (N11001, N10941_t1, N8655);
not NOT1_3324 (N11002, N10944_t0);
nand NAND2_3325 (N11003, N10944_t1, N9456);
not NOT1_3326 (N11004, N10947_t0);
nand NAND2_3327 (N11005, N10947_t1, N9461);
not NOT1_3328 (N11006, N10950_t0);
nand NAND2_3329 (N11007, N10950_t1, N9465);
nand NAND2_3330 (N11008, N10981, N10954);
not NOT1_3331 (N11011, N10955_t0);
nand NAND2_3332 (N11012, N10955_t1, N9495);
not NOT1_3333 (N11013, N10958_t0);
nand NAND2_3334 (N11014, N10958_t1, N9500);
nand NAND2_3335 (N11015, N10986, N10962);
nand NAND2_3336 (N11018, N10987, N10964);
nand NAND2_3337 (N11023, N7453_t1, N10988);
nand NAND2_3338 (N11024, N7471_t1, N10990);
nand NAND2_3339 (N11027, N7509_t1, N10998);
nand NAND2_3340 (N11028, N7527_t1, N11000);
nand NAND2_3341 (N11029, N8684_t1, N11002);
nand NAND2_3342 (N11030, N8696_t1, N11004);
nand NAND2_3343 (N11031, N8702_t1, N11006);
nand NAND2_3344 (N11034, N8763_t1, N11011);
nand NAND2_3345 (N11035, N8775_t1, N11013);
not NOT1_3346 (N11040, N10992_t0);
nand NAND2_3347 (N11041, N10992_t1, N8294);
not NOT1_3348 (N11042, N10995_t0);
nand NAND2_3349 (N11043, N10995_t1, N8295);
nand NAND2_3350 (N11044, N11023, N10989);
nand NAND2_3351 (N11047, N11024, N10991);
nand NAND2_3352 (N11050, N11027, N10999);
nand NAND2_3353 (N11053, N11028, N11001);
nand NAND2_3354 (N11056, N11029, N11003);
nand NAND2_3355 (N11059, N11030, N11005);
nand NAND2_3356 (N11062, N11031, N11007);
not NOT1_3357 (N11065, N11008_t0);
nand NAND2_3358 (N11066, N11008_t1, N9477);
nand NAND2_3359 (N11067, N11034, N11012);
nand NAND2_3360 (N11070, N11035, N11014);
not NOT1_3361 (N11073, N11015_t0);
nand NAND2_3362 (N11074, N11015_t1, N9507);
not NOT1_3363 (N11075, N11018_t0);
nand NAND2_3364 (N11076, N11018_t1, N9516);
nand NAND2_3365 (N11077, N7488_t1, N11040);
nand NAND2_3366 (N11078, N7500_t1, N11042);
nand NAND2_3367 (N11095, N8721_t1, N11065);
nand NAND2_3368 (N11098, N8787_t1, N11073);
nand NAND2_3369 (N11099, N8805_t1, N11075);
nand NAND2_3370 (N11100, N11077, N11041);
nand NAND2_3371 (N11103, N11078, N11043);
not NOT1_3372 (N11106, N11056_t0);
nand NAND2_3373 (N11107, N11056_t1, N9319);
not NOT1_3374 (N11108, N11059_t0);
nand NAND2_3375 (N11109, N11059_t1, N9320);
not NOT1_3376 (N11110, N11067_t0);
nand NAND2_3377 (N11111, N11067_t1, N9381);
not NOT1_3378 (N11112, N11070_t0);
nand NAND2_3379 (N11113, N11070_t1, N9382);
not NOT1_3380 (N11114, N11044_t0);
nand NAND2_3381 (N11115, N11044_t1, N8618);
not NOT1_3382 (N11116, N11047_t0);
nand NAND2_3383 (N11117, N11047_t1, N8619);
not NOT1_3384 (N11118, N11050_t0);
nand NAND2_3385 (N11119, N11050_t1, N8647);
not NOT1_3386 (N11120, N11053_t0);
nand NAND2_3387 (N11121, N11053_t1, N8648);
not NOT1_3388 (N11122, N11062_t0);
nand NAND2_3389 (N11123, N11062_t1, N9466);
nand NAND2_3390 (N11124, N11095, N11066);
nand NAND2_3391 (N11127, N11098, N11074);
nand NAND2_3392 (N11130, N11099, N11076);
nand NAND2_3393 (N11137, N8687_t1, N11106);
nand NAND2_3394 (N11138, N8699_t1, N11108);
nand NAND2_3395 (N11139, N8766_t1, N11110);
nand NAND2_3396 (N11140, N8778_t1, N11112);
nand NAND2_3397 (N11141, N7456_t1, N11114);
nand NAND2_3398 (N11142, N7474_t1, N11116);
nand NAND2_3399 (N11143, N7512_t1, N11118);
nand NAND2_3400 (N11144, N7530_t1, N11120);
nand NAND2_3401 (N11145, N8705_t1, N11122);
and AND3_3402 (N11152, N11103_t0, N8871_t1, N10283_t0);
and AND3_3403 (N11153, N11100_t0, N7655_t2, N10283_t1);
and AND3_3404 (N11154, N11103_t1, N9551_t1, N10119_t1);
and AND3_3405 (N11155, N11100_t1, N9917, N10119_t2);
nand NAND2_3406 (N11156, N11137, N11107);
nand NAND2_3407 (N11159, N11138, N11109);
nand NAND2_3408 (N11162, N11139, N11111);
nand NAND2_3409 (N11165, N11140, N11113);
nand NAND2_3410 (N11168, N11141, N11115);
nand NAND2_3411 (N11171, N11142, N11117);
nand NAND2_3412 (N11174, N11143, N11119);
nand NAND2_3413 (N11177, N11144, N11121);
nand NAND2_3414 (N11180, N11145, N11123);
not NOT1_3415 (N11183, N11124_t0);
nand NAND2_3416 (N11184, N11124_t1, N9468);
not NOT1_3417 (N11185, N11127_t0);
nand NAND2_3418 (N11186, N11127_t1, N9508);
not NOT1_3419 (N11187, N11130_t0);
nand NAND2_3420 (N11188, N11130_t1, N9509);
or OR4_3421 (N11205, N11152, N11153, N11154, N11155);
nand NAND2_3422 (N11210, N8724_t1, N11183);
nand NAND2_3423 (N11211, N8790_t1, N11185);
nand NAND2_3424 (N11212, N8808_t1, N11187);
not NOT1_3425 (N11213, N11168_t0);
nand NAND2_3426 (N11214, N11168_t1, N8260);
not NOT1_3427 (N11215, N11171_t0);
nand NAND2_3428 (N11216, N11171_t1, N8261);
not NOT1_3429 (N11217, N11174_t0);
nand NAND2_3430 (N11218, N11174_t1, N8296);
not NOT1_3431 (N11219, N11177_t0);
nand NAND2_3432 (N11220, N11177_t1, N8297);
and AND3_3433 (N11222, N11159_t0, N9575_t2, N1218_t0);
and AND3_3434 (N11223, N11156_t0, N8927_t2, N1218_t1);
and AND3_3435 (N11224, N11159_t1, N9935_t1, N750_t1);
and AND3_3436 (N11225, N11156_t1, N10132, N750_t2);
and AND3_3437 (N11226, N11165_t0, N9608_t1, N10497_t0);
and AND3_3438 (N11227, N11162_t0, N9001_t2, N10497_t1);
and AND3_3439 (N11228, N11165_t1, N9949_t1, N10301_t1);
and AND3_3440 (N11229, N11162_t1, N10160, N10301_t2);
not NOT1_3441 (N11231, N11180_t0);
nand NAND2_3442 (N11232, N11180_t1, N9467);
nand NAND2_3443 (N11233, N11210, N11184);
nand NAND2_3444 (N11236, N11211, N11186);
nand NAND2_3445 (N11239, N11212, N11188);
nand NAND2_3446 (N11242, N7459_t1, N11213);
nand NAND2_3447 (N11243, N7462_t1, N11215);
nand NAND2_3448 (N11244, N7515_t1, N11217);
nand NAND2_3449 (N11245, N7518_t1, N11219);
not NOT1_3450 (N11246, N11205_t0);
nand NAND2_3451 (N11250, N8708_t1, N11231);
or OR4_3452 (N11252, N11222, N11223, N11224, N11225);
or OR4_3453 (N11257, N11226, N11227, N11228, N11229);
nand NAND2_3454 (N11260, N11242, N11214);
nand NAND2_3455 (N11261, N11243, N11216);
nand NAND2_3456 (N11262, N11244, N11218);
nand NAND2_3457 (N11263, N11245, N11220);
not NOT1_3458 (N11264, N11233_t0);
nand NAND2_3459 (N11265, N11233_t1, N9322);
not NOT1_3460 (N11267, N11236_t0);
nand NAND2_3461 (N11268, N11236_t1, N9383);
not NOT1_3462 (N11269, N11239_t0);
nand NAND2_3463 (N11270, N11239_t1, N9384);
nand NAND2_3464 (N11272, N11250, N11232);
not NOT1_3465 (N11277, N11261);
and AND2_3466 (N11278, N10273_t3, N11260);
not NOT1_3467 (N11279, N11263);
and AND2_3468 (N11280, N10119_t3, N11262);
nand NAND2_3469 (N11282, N8714_t1, N11264);
not NOT1_3470 (N11283, N11252_t0);
nand NAND2_3471 (N11284, N8793_t1, N11267);
nand NAND2_3472 (N11285, N8796_t1, N11269);
not NOT1_3473 (N11286, N11257_t0);
and AND2_3474 (N11288, N11277, N10479_t2);
and AND2_3475 (N11289, N11279, N10283_t2);
not NOT1_3476 (N11290, N11272_t0);
nand NAND2_3477 (N11291, N11272_t1, N9321);
nand NAND2_3478 (N11292, N11282, N11265);
nand NAND2_3479 (N11293, N11284, N11268);
nand NAND2_3480 (N11294, N11285, N11270);
nand NAND2_3481 (N11295, N8711_t1, N11290);
not NOT1_3482 (N11296, N11292);
not NOT1_3483 (N11297, N11294);
and AND2_3484 (N11298, N10301_t3, N11293);
or OR2_3485 (N11299, N11288, N11278);
or OR2_3486 (N11302, N11289, N11280);
nand NAND2_3487 (N11307, N11295, N11291);
and AND2_3488 (N11308, N11296, N1218_t2);
and AND2_3489 (N11309, N11297, N10497_t2);
nand NAND2_3490 (N11312, N11302_t0, N11246);
nand NAND2_3491 (N11313, N11299_t0, N10836);
not NOT1_3492 (N11314, N11299_t1);
not NOT1_3493 (N11315, N11302_t1);
and AND2_3494 (N11316, N750_t3, N11307);
or OR2_3495 (N11317, N11309, N11298);
nand NAND2_3496 (N11320, N11205_t1, N11315);
nand NAND2_3497 (N11321, N10739_t1, N11314);
or OR2_3498 (N11323, N11308, N11316);
nand NAND2_3499 (N11327, N11312, N11320);
nand NAND2_3500 (N11328, N11313, N11321);
nand NAND2_3501 (N11329, N11317_t0, N11286);
not NOT1_3502 (N11331, N11317_t1);
not NOT1_3503 (N11333, N11327);
not NOT1_3504 (N11334, N11328);
nand NAND2_3505 (N11335, N11257_t1, N11331);
nand NAND2_3506 (N11336, N11323_t0, N11283);
not NOT1_3507 (N11337, N11323_t1);
nand NAND2_3508 (N11338, N11329, N11335);
nand NAND2_3509 (N11339, N11252_t1, N11337);
not NOT1_3510 (N11340, N11338);
nand NAND2_3511 (N11341, N11336, N11339);
not NOT1_3512 (N11342, N11341);
buf BUFF1_3513 (N241_O, N241_I_t);

endmodule
