/* 
    Fault Injection Circuitry

    Injects Faults in CUT
*/

module fic (
);
    
endmodule