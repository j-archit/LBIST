/* 
    Test Pattern Generator

    Consists of 
    1. Random Pattern Generator (rpg.v)
    2. Deterministic Pattern Generator (dpg.v)
    3. Selection Multiplexer

*/

module tpg
#(parameter INPUT_BITS = 4)
(
    input type
);
    
endmodule