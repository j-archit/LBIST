// Verilog
// c3540
// Ninputs 50
// Noutputs 22
// NtotalGates 1669
// BUFF1 223
// NOT1 490
// OR2 35
// AND2 410
// NAND2 274
// NAND3 17
// AND3 76
// NOR2 25
// AND4 10
// NAND4 7
// OR3 56
// NOR3 27
// AND5 2
// NOR8 16
// OR4 1

module c3540f (INC,END,clk,rst,N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
              N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
              N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
              N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
              N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,
              N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
              N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
              N5360,N5361);

input N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
      N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
      N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
      N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
      N303,N311,N317,N322,N326,N329,N330,N343,N349,N350;

output N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
       N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
       N5360,N5361;

wire N655,N665,N670,N679,N683,N686,N690,N699,N702,N706,
     N715,N724,N727,N736,N740,N749,N753,N763,N768,N769,
     N772,N779,N782,N786,N793,N794,N798,N803,N820,N821,
     N825,N829,N832,N835,N836,N839,N842,N845,N848,N851,
     N854,N858,N861,N864,N867,N870,N874,N877,N880,N883,
     N886,N889,N890,N891,N892,N895,N896,N913,N914,N915,
     N916,N917,N920,N923,N926,N929,N932,N935,N938,N941,
     N944,N947,N950,N953,N956,N959,N962,N965,N1067,N1117,
     N1179,N1196,N1197,N1202,N1219,N1250,N1251,N1252,N1253,N1254,
     N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
     N1267,N1268,N1271,N1272,N1273,N1276,N1279,N1298,N1302,N1306,
     N1315,N1322,N1325,N1328,N1331,N1334,N1337,N1338,N1339,N1340,
     N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
     N1353,N1358,N1363,N1366,N1369,N1384,N1401,N1402,N1403,N1404,
     N1405,N1406,N1407,N1408,N1409,N1426,N1427,N1452,N1459,N1460,
     N1461,N1464,N1467,N1468,N1469,N1470,N1471,N1474,N1475,N1478,
     N1481,N1484,N1487,N1490,N1493,N1496,N1499,N1502,N1505,N1507,
     N1508,N1509,N1510,N1511,N1512,N1520,N1562,N1579,N1580,N1581,
     N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,
     N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1643,
     N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1667,N1670,N1673,
     N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1691,N1692,N1693,
     N1694,N1714,N1715,N1718,N1721,N1722,N1725,N1726,N1727,N1728,
     N1729,N1730,N1731,N1735,N1736,N1737,N1738,N1747,N1756,N1761,
     N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1787,N1788,N1789,
     N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,
     N1800,N1801,N1802,N1803,N1806,N1809,N1812,N1815,N1818,N1821,
     N1824,N1833,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
     N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
     N1860,N1861,N1862,N1863,N1864,N1869,N1870,N1873,N1874,N1875,
     N1878,N1879,N1880,N1883,N1884,N1885,N1888,N1889,N1890,N1893,
     N1894,N1895,N1898,N1899,N1900,N1903,N1904,N1905,N1908,N1909,
     N1912,N1913,N1917,N1922,N1926,N1930,N1933,N1936,N1939,N1940,
     N1941,N1942,N1943,N1944,N1945,N1946,N1960,N1961,N1966,N1981,
     N1982,N1983,N1986,N1987,N1988,N1989,N1990,N1991,N2022,N2023,
     N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
     N2034,N2035,N2036,N2037,N2038,N2043,N2052,N2057,N2068,N2073,
     N2078,N2083,N2088,N2093,N2098,N2103,N2121,N2122,N2123,N2124,
     N2125,N2126,N2127,N2128,N2133,N2134,N2135,N2136,N2137,N2138,
     N2139,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,
     N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2175,
     N2178,N2179,N2180,N2181,N2183,N2184,N2185,N2188,N2191,N2194,
     N2197,N2200,N2203,N2206,N2209,N2210,N2211,N2212,N2221,N2230,
     N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,
     N2241,N2242,N2243,N2244,N2245,N2270,N2277,N2282,N2287,N2294,
     N2299,N2304,N2307,N2310,N2313,N2316,N2319,N2322,N2325,N2328,
     N2331,N2334,N2341,N2342,N2347,N2348,N2349,N2350,N2351,N2352,
     N2353,N2354,N2355,N2374,N2375,N2376,N2379,N2398,N2417,N2418,
     N2419,N2420,N2421,N2422,N2425,N2426,N2427,N2430,N2431,N2432,
     N2435,N2436,N2437,N2438,N2439,N2440,N2443,N2444,N2445,N2448,
     N2449,N2450,N2467,N2468,N2469,N2470,N2471,N2474,N2475,N2476,
     N2477,N2478,N2481,N2482,N2483,N2486,N2487,N2488,N2497,N2506,
     N2515,N2524,N2533,N2542,N2551,N2560,N2569,N2578,N2587,N2596,
     N2605,N2614,N2623,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
     N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,
     N2652,N2656,N2659,N2662,N2666,N2670,N2673,N2677,N2681,N2684,
     N2688,N2692,N2697,N2702,N2706,N2710,N2715,N2719,N2723,N2728,
     N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
     N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2748,N2749,
     N2750,N2751,N2754,N2755,N2756,N2757,N2758,N2761,N2764,N2768,
     N2769,N2898,N2899,N2900,N2901,N2962,N2966,N2967,N2970,N2973,
     N2977,N2980,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,
     N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
     N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,
     N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,
     N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,
     N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,
     N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,
     N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,
     N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,
     N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,
     N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,
     N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,
     N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,
     N3112,N3115,N3118,N3119,N3122,N3125,N3128,N3131,N3134,N3135,
     N3138,N3141,N3142,N3145,N3148,N3149,N3152,N3155,N3158,N3161,
     N3164,N3165,N3168,N3171,N3172,N3175,N3178,N3181,N3184,N3187,
     N3190,N3191,N3192,N3193,N3194,N3196,N3206,N3207,N3208,N3209,
     N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,
     N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,
     N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,
     N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,
     N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,
     N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,
     N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,
     N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,
     N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,
     N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,
     N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,
     N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,
     N3330,N3331,N3332,N3333,N3334,N3383,N3384,N3387,N3388,N3389,
     N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,
     N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3410,N3413,
     N3414,N3415,N3419,N3423,N3426,N3429,N3430,N3431,N3434,N3437,
     N3438,N3439,N3442,N3445,N3446,N3447,N3451,N3455,N3458,N3461,
     N3462,N3463,N3466,N3469,N3470,N3471,N3472,N3475,N3478,N3481,
     N3484,N3487,N3490,N3493,N3496,N3499,N3502,N3505,N3508,N3511,
     N3514,N3517,N3520,N3523,N3534,N3535,N3536,N3537,N3538,N3539,
     N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,
     N3550,N3551,N3552,N3557,N3568,N3573,N3578,N3589,N3594,N3605,
     N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,
     N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
     N3648,N3651,N3652,N3653,N3654,N3657,N3658,N3661,N3662,N3663,
     N3664,N3667,N3670,N3671,N3672,N3673,N3676,N3677,N3680,N3681,
     N3682,N3685,N3686,N3687,N3688,N3689,N3690,N3693,N3694,N3695,
     N3696,N3697,N3700,N3703,N3704,N3705,N3706,N3707,N3708,N3711,
     N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,
     N3731,N3734,N3740,N3743,N3753,N3756,N3762,N3765,N3766,N3773,
     N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3786,N3789,N3800,
     N3803,N3809,N3812,N3815,N3818,N3821,N3824,N3827,N3830,N3834,
     N3835,N3838,N3845,N3850,N3855,N3858,N3861,N3865,N3868,N3884,
     N3885,N3894,N3895,N3898,N3899,N3906,N3911,N3912,N3913,N3916,
     N3917,N3920,N3921,N3924,N3925,N3926,N3930,N3931,N3932,N3935,
     N3936,N3937,N3940,N3947,N3948,N3950,N3953,N3956,N3959,N3962,
     N3965,N3968,N3971,N3974,N3977,N3980,N3983,N3992,N3996,N4013,
     N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4042,N4043,N4044,
     N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,
     N4055,N4056,N4057,N4058,N4059,N4062,N4065,N4066,N4067,N4070,
     N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4085,N4086,
     N4088,N4090,N4091,N4094,N4098,N4101,N4104,N4105,N4106,N4107,
     N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4119,
     N4122,N4123,N4126,N4127,N4128,N4139,N4142,N4146,N4147,N4148,
     N4149,N4150,N4151,N4152,N4153,N4154,N4161,N4167,N4174,N4182,
     N4186,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
     N4200,N4203,N4209,N4213,N4218,N4223,N4238,N4239,N4241,N4242,
     N4247,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4283,
     N4284,N4287,N4291,N4295,N4296,N4299,N4303,N4304,N4305,N4310,
     N4316,N4317,N4318,N4319,N4322,N4325,N4326,N4327,N4328,N4329,
     N4330,N4331,N4335,N4338,N4341,N4344,N4347,N4350,N4353,N4356,
     N4359,N4362,N4365,N4368,N4371,N4376,N4377,N4387,N4390,N4393,
     N4398,N4413,N4416,N4421,N4427,N4430,N4435,N4442,N4443,N4446,
     N4447,N4448,N4452,N4458,N4461,N4462,N4463,N4464,N4465,N4468,
     N4472,N4475,N4479,N4484,N4486,N4487,N4491,N4493,N4496,N4497,
     N4498,N4503,N4506,N4507,N4508,N4509,N4510,N4511,N4515,N4526,
     N4527,N4528,N4529,N4530,N4531,N4534,N4537,N4540,N4545,N4549,
     N4552,N4555,N4558,N4559,N4562,N4563,N4564,N4568,N4569,N4572,
     N4573,N4576,N4581,N4584,N4587,N4588,N4593,N4596,N4597,N4599,
     N4602,N4603,N4608,N4613,N4616,N4619,N4623,N4628,N4629,N4630,
     N4635,N4636,N4640,N4641,N4642,N4643,N4644,N4647,N4650,N4656,
     N4659,N4664,N4668,N4669,N4670,N4673,N4674,N4675,N4676,N4677,
     N4678,N4679,N4687,N4688,N4691,N4694,N4697,N4700,N4704,N4705,
     N4706,N4707,N4708,N4711,N4716,N4717,N4721,N4722,N4726,N4727,
     N4730,N4733,N4740,N4743,N4747,N4748,N4749,N4750,N4753,N4754,
     N4755,N4756,N4757,N4769,N4772,N4775,N4778,N4786,N4787,N4788,
     N4789,N4794,N4797,N4800,N4805,N4808,N4812,N4816,N4817,N4818,
     N4822,N4823,N4826,N4829,N4830,N4831,N4838,N4844,N4847,N4850,
     N4854,N4859,N4860,N4868,N4870,N4872,N4873,N4876,N4880,N4885,
     N4889,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4904,
     N4905,N4906,N4907,N4913,N4916,N4920,N4921,N4924,N4925,N4926,
     N4928,N4929,N4930,N4931,N4937,N4940,N4946,N4949,N4950,N4951,
     N4952,N4953,N4954,N4957,N4964,N4965,N4968,N4969,N4970,N4973,
     N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4988,N4991,
     N4996,N4999,N5007,N5010,N5013,N5018,N5021,N5026,N5029,N5030,
     N5039,N5042,N5046,N5050,N5055,N5058,N5061,N5066,N5070,N5080,
     N5085,N5094,N5095,N5097,N5103,N5108,N5109,N5110,N5111,N5114,
     N5117,N5122,N5125,N5128,N5133,N5136,N5139,N5145,N5151,N5154,
     N5159,N5160,N5163,N5166,N5173,N5174,N5177,N5182,N5183,N5184,
     N5188,N5193,N5196,N5197,N5198,N5199,N5201,N5203,N5205,N5209,
     N5212,N5215,N5217,N5219,N5220,N5221,N5222,N5223,N5224,N5225,
     N5228,N5232,N5233,N5234,N5235,N5236,N5240,N5242,N5243,N5245,
     N5246,N5250,N5253,N5254,N5257,N5258,N5261,N5266,N5269,N5277,
     N5278,N5279,N5283,N5284,N5285,N5286,N5289,N5292,N5295,N5298,
     N5303,N5306,N5309,N5312,N5313,N5322,N5323,N5324,N5327,N5332,
     N5335,N5340,N5341,N5344,N5345,N5348,N5349,N5350,N5351,N5352,
     N5353,N5354,N5355,N5356,N5357,N5358,N5359;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N124_t,N222_t,N329_t,N349_t;
wire N50_t0,N50_t1,N50_t2,N50_t3,N50_t4,N50_t5,N50_t6,N58_t0,N58_t1,
     N58_t2,N58_t3,N58_t4,N58_t5,N58_t6,N58_t7,N58_t8,N68_t0,N68_t1,N68_t2,
     N68_t3,N68_t4,N68_t5,N68_t6,N68_t7,N77_t0,N77_t1,N77_t2,N77_t3,N77_t4,
     N77_t5,N77_t6,N77_t7,N77_t8,N87_t0,N87_t1,N87_t2,N87_t3,N87_t4,N87_t5,
     N87_t6,N87_t7,N87_t8,N97_t0,N97_t1,N97_t2,N97_t3,N97_t4,N97_t5,N97_t6,
     N97_t7,N97_t8,N107_t0,N107_t1,N107_t2,N107_t3,N107_t4,N107_t5,N107_t6,N107_t7,
     N116_t0,N116_t1,N116_t2,N116_t3,N116_t4,N116_t5,N116_t6,N257_t0,N257_t1,N257_t2,
     N257_t3,N257_t4,N257_t5,N264_t0,N264_t1,N264_t2,N264_t3,N264_t4,N1_t0,N1_t1,
     N1_t2,N1_t3,N1_t4,N1_t5,N1_t6,N1_t7,N1_t8,N1_t9,N1_t10,N13_t0,
     N13_t1,N13_t2,N13_t3,N13_t4,N13_t5,N20_t0,N20_t1,N20_t2,N20_t3,N20_t4,
     N20_t5,N20_t6,N20_t7,N20_t8,N20_t9,N20_t10,N20_t11,N33_t0,N33_t1,N33_t2,
     N33_t3,N33_t4,N33_t5,N33_t6,N41_t0,N41_t1,N41_t2,N45_t0,N45_t1,N45_t2,
     N45_t3,N190_t0,N190_t1,N190_t2,N190_t3,N190_t4,N190_t5,N190_t6,N190_t7,N190_t8,
     N200_t0,N200_t1,N200_t2,N200_t3,N200_t4,N200_t5,N200_t6,N200_t7,N200_t8,N200_t9,
     N200_t10,N200_t11,N179_t0,N179_t1,N179_t2,N179_t3,N179_t4,N179_t5,N179_t6,N179_t7,
     N179_t8,N179_t9,N213_t0,N213_t1,N213_t2,N213_t3,N213_t4,N213_t5,N213_t6,N213_t7,
     N343_t0,N343_t1,N343_t2,N343_t3,N343_t4,N226_t0,N226_t1,N226_t2,N226_t3,N226_t4,
     N232_t0,N232_t1,N232_t2,N232_t3,N232_t4,N238_t0,N238_t1,N238_t2,N238_t3,N238_t4,
     N244_t0,N244_t1,N244_t2,N244_t3,N244_t4,N250_t0,N250_t1,N250_t2,N250_t3,N250_t4,
     N250_t5,N270_t0,N270_t1,N270_t2,N330_t0,N330_t1,N330_t2,N330_t3,N330_t4,N330_t5,
     N330_t6,N330_t7,N330_t8,N330_t9,N330_t10,N330_t11,N169_t0,N169_t1,N169_t2,N169_t3,
     N169_t4,N169_t5,N169_t6,N169_t7,N169_t8,N842_t0,N842_t1,N848_t0,N848_t1,N854_t0,
     N854_t1,N854_t2,N655_t0,N655_t1,N655_t2,N655_t3,N655_t4,N655_t5,N655_t6,N655_t7,
     N655_t8,N670_t0,N670_t1,N670_t2,N670_t3,N670_t4,N670_t5,N670_t6,N670_t7,N690_t0,
     N690_t1,N690_t2,N690_t3,N690_t4,N690_t5,N690_t6,N690_t7,N706_t0,N706_t1,N706_t2,
     N706_t3,N706_t4,N706_t5,N706_t6,N706_t7,N715_t0,N715_t1,N715_t2,N715_t3,N715_t4,
     N715_t5,N715_t6,N715_t7,N727_t0,N727_t1,N727_t2,N727_t3,N727_t4,N727_t5,N727_t6,
     N727_t7,N740_t0,N740_t1,N740_t2,N740_t3,N740_t4,N740_t5,N740_t6,N740_t7,N753_t0,
     N753_t1,N753_t2,N753_t3,N753_t4,N753_t5,N753_t6,N753_t7,N753_t8,N926_t0,N926_t1,
     N929_t0,N929_t1,N932_t0,N932_t1,N935_t0,N935_t1,N679_t0,N679_t1,N679_t2,N686_t0,
     N686_t1,N686_t2,N736_t0,N736_t1,N736_t2,N749_t0,N749_t1,N749_t2,N683_t0,N683_t1,
     N699_t0,N699_t1,N665_t0,N665_t1,N665_t2,N665_t3,N953_t0,N953_t1,N959_t0,N959_t1,
     N839_t0,N839_t1,N782_t0,N782_t1,N782_t2,N825_t0,N825_t1,N825_t2,N832_t0,N832_t1,
     N779_t0,N779_t1,N836_t0,N836_t1,N769_t0,N769_t1,N772_t0,N772_t1,N772_t2,N772_t3,
     N772_t4,N772_t5,N786_t0,N786_t1,N786_t2,N786_t3,N786_t4,N786_t5,N798_t0,N798_t1,
     N798_t2,N798_t3,N874_t0,N874_t1,N794_t0,N794_t1,N794_t2,N956_t0,N956_t1,N861_t0,
     N861_t1,N867_t0,N867_t1,N870_t0,N870_t1,N870_t2,N962_t0,N962_t1,N803_t0,N803_t1,
     N803_t2,N803_t3,N803_t4,N803_t5,N803_t6,N803_t7,N803_t8,N803_t9,N803_t10,N803_t11,
     N803_t12,N803_t13,N803_t14,N803_t15,N883_t0,N883_t1,N886_t0,N886_t1,N892_t0,N892_t1,
     N821_t0,N821_t1,N821_t2,N896_t0,N896_t1,N896_t2,N896_t3,N896_t4,N896_t5,N896_t6,
     N896_t7,N896_t8,N896_t9,N896_t10,N896_t11,N896_t12,N896_t13,N896_t14,N896_t15,N829_t0,
     N829_t1,N917_t0,N917_t1,N965_t0,N965_t1,N920_t0,N920_t1,N923_t0,N923_t1,N938_t0,
     N938_t1,N941_t0,N941_t1,N944_t0,N944_t1,N947_t0,N947_t1,N950_t0,N950_t1,N702_t0,
     N702_t1,N702_t2,N724_t0,N724_t1,N763_t0,N763_t1,N763_t2,N763_t3,N877_t0,N877_t1,
     N880_t0,N880_t1,N1117_t0,N1117_t1,N1117_t2,N1117_t3,N1117_t4,N1117_t5,N1117_t6,N1117_t7,
     N1117_t8,N1117_t9,N1117_t10,N1117_t11,N1117_t12,N1117_t13,N1117_t14,N1117_t15,N223_t0,N223_t1,
     N1202_t0,N1202_t1,N1202_t2,N1202_t3,N1202_t4,N1202_t5,N1202_t6,N1202_t7,N1202_t8,N1202_t9,
     N1202_t10,N1202_t11,N1202_t12,N1202_t13,N1202_t14,N1202_t15,N1264_t0,N1264_t1,N1340_t0,N1340_t1,
     N1268_t0,N1268_t1,N1493_t0,N1493_t1,N1499_t0,N1499_t1,N1273_t0,N1273_t1,N1276_t0,N1276_t1,
     N1325_t0,N1325_t1,N1279_t0,N1279_t1,N1302_t0,N1302_t1,N1302_t2,N1496_t0,N1496_t1,N1502_t0,
     N1502_t1,N1328_t0,N1328_t1,N1334_t0,N1334_t1,N1331_t0,N1331_t1,N845_t0,N845_t1,N150_t0,
     N150_t1,N150_t2,N150_t3,N150_t4,N150_t5,N150_t6,N150_t7,N851_t0,N851_t1,N159_t0,
     N159_t1,N159_t2,N159_t3,N159_t4,N159_t5,N159_t6,N159_t7,N159_t8,N858_t0,N858_t1,
     N864_t0,N864_t1,N283_t0,N283_t1,N283_t2,N283_t3,N283_t4,N283_t5,N283_t6,N283_t7,
     N283_t8,N283_t9,N1363_t0,N1363_t1,N1366_t0,N1366_t1,N1298_t0,N1298_t1,N1298_t2,N1369_t0,
     N1369_t1,N1369_t2,N1369_t3,N1369_t4,N1369_t5,N1369_t6,N1369_t7,N1369_t8,N1369_t9,N1369_t10,
     N1369_t11,N1369_t12,N1369_t13,N1384_t0,N1384_t1,N1384_t2,N1384_t3,N1384_t4,N1384_t5,N1384_t6,
     N1384_t7,N1384_t8,N1384_t9,N1384_t10,N1384_t11,N1384_t12,N1384_t13,N1384_t14,N1384_t15,N1409_t0,
     N1409_t1,N1409_t2,N1409_t3,N1409_t4,N1409_t5,N1409_t6,N1409_t7,N1409_t8,N1409_t9,N1409_t10,
     N1409_t11,N1409_t12,N1409_t13,N1409_t14,N1409_t15,N1306_t0,N1306_t1,N1306_t2,N1306_t3,N1306_t4,
     N1306_t5,N1306_t6,N1306_t7,N1322_t0,N1322_t1,N1315_t0,N1315_t1,N1315_t2,N1315_t3,N1315_t4,
     N1315_t5,N1452_t0,N1452_t1,N1452_t2,N1452_t3,N1452_t4,N1452_t5,N1464_t0,N1464_t1,N1471_t0,
     N1471_t1,N1475_t0,N1475_t1,N1478_t0,N1478_t1,N1481_t0,N1481_t1,N1484_t0,N1484_t1,N1487_t0,
     N1487_t1,N1490_t0,N1490_t1,N1520_t0,N1520_t1,N1520_t2,N294_t0,N294_t1,N294_t2,N294_t3,
     N294_t4,N294_t5,N294_t6,N294_t7,N303_t0,N303_t1,N303_t2,N303_t3,N303_t4,N303_t5,
     N303_t6,N1667_t0,N1667_t1,N1670_t0,N1670_t1,N1197_t0,N1197_t1,N1197_t2,N1197_t3,N1219_t0,
     N1219_t1,N1219_t2,N1219_t3,N1562_t0,N1562_t1,N1562_t2,N1562_t3,N1562_t4,N1562_t5,N1562_t6,
     N1562_t7,N1562_t8,N1562_t9,N1562_t10,N1562_t11,N1562_t12,N1562_t13,N1562_t14,N1562_t15,N1933_t0,
     N1933_t1,N1936_t0,N1936_t1,N1738_t0,N1738_t1,N1738_t2,N1738_t3,N1738_t4,N1738_t5,N1738_t6,
     N1738_t7,N1747_t0,N1747_t1,N1747_t2,N1747_t3,N1747_t4,N1747_t5,N1747_t6,N1747_t7,N1722_t0,
     N1722_t1,N1761_t0,N1761_t1,N1756_t0,N1756_t1,N1756_t2,N1756_t3,N1358_t0,N1358_t1,N1358_t2,
     N1358_t3,N1812_t0,N1812_t1,N1809_t0,N1809_t1,N1353_t0,N1353_t1,N1353_t2,N1353_t3,N1806_t0,
     N1806_t1,N1803_t0,N1803_t1,N1815_t0,N1815_t1,N1818_t0,N1818_t1,N1821_t0,N1821_t1,N1833_t0,
     N1833_t1,N1833_t2,N1833_t3,N1833_t4,N1833_t5,N1833_t6,N1833_t7,N1824_t0,N1824_t1,N1824_t2,
     N1824_t3,N1824_t4,N1824_t5,N1824_t6,N1824_t7,N1917_t0,N1917_t1,N1917_t2,N1917_t3,N1930_t0,
     N1930_t1,N350_t0,N350_t1,N1715_t0,N1715_t1,N1718_t0,N1718_t1,N2057_t0,N2057_t1,N2057_t2,
     N2057_t3,N2057_t4,N2057_t5,N2057_t6,N2057_t7,N274_t0,N274_t1,N274_t2,N274_t3,N274_t4,
     N274_t5,N274_t6,N274_t7,N2052_t0,N2052_t1,N2052_t2,N2052_t3,N2043_t0,N2043_t1,N2043_t2,
     N2043_t3,N2043_t4,N2043_t5,N2043_t6,N2043_t7,N2038_t0,N2038_t1,N2038_t2,N2038_t3,N2313_t0,
     N2313_t1,N2316_t0,N2316_t1,N2319_t0,N2319_t1,N2322_t0,N2322_t1,N2325_t0,N2325_t1,N2328_t0,
     N2328_t1,N2331_t0,N2331_t1,N2334_t0,N2334_t1,N2175_t0,N2175_t1,N2185_t0,N2185_t1,N2188_t0,
     N2188_t1,N2191_t0,N2191_t1,N2194_t0,N2194_t1,N2197_t0,N2197_t1,N2200_t0,N2200_t1,N2203_t0,
     N2203_t1,N2206_t0,N2206_t1,N2212_t0,N2212_t1,N2212_t2,N2212_t3,N2212_t4,N2212_t5,N2212_t6,
     N2212_t7,N2221_t0,N2221_t1,N2221_t2,N2221_t3,N2221_t4,N2221_t5,N2221_t6,N2221_t7,N2270_t0,
     N2270_t1,N1870_t0,N1870_t1,N2068_t0,N2068_t1,N2277_t0,N2277_t1,N1880_t0,N1880_t1,N2078_t0,
     N2078_t1,N2282_t0,N2282_t1,N1885_t0,N1885_t1,N2083_t0,N2083_t1,N2287_t0,N2287_t1,N1890_t0,
     N1890_t1,N2088_t0,N2088_t1,N2294_t0,N2294_t1,N1900_t0,N1900_t1,N2098_t0,N2098_t1,N2299_t0,
     N2299_t1,N1905_t0,N1905_t1,N2103_t0,N2103_t1,N2304_t0,N2304_t1,N2158_t0,N2158_t1,N2158_t2,
     N2158_t3,N2158_t4,N2158_t5,N2158_t6,N2158_t7,N2158_t8,N2158_t9,N2158_t10,N2158_t11,N2158_t12,
     N2158_t13,N2158_t14,N2158_t15,N2376_t0,N2376_t1,N1983_t0,N1983_t1,N2379_t0,N2379_t1,N2471_t0,
     N2471_t1,N2488_t0,N2488_t1,N2488_t2,N2488_t3,N2488_t4,N2488_t5,N2488_t6,N2488_t7,N2497_t0,
     N2497_t1,N2497_t2,N2497_t3,N2497_t4,N2497_t5,N2497_t6,N2497_t7,N2506_t0,N2506_t1,N2506_t2,
     N2506_t3,N2506_t4,N2506_t5,N2506_t6,N2506_t7,N2515_t0,N2515_t1,N2515_t2,N2515_t3,N2515_t4,
     N2515_t5,N2515_t6,N2515_t7,N2524_t0,N2524_t1,N2524_t2,N2524_t3,N2524_t4,N2524_t5,N2524_t6,
     N2524_t7,N2533_t0,N2533_t1,N2533_t2,N2533_t3,N2533_t4,N2533_t5,N2533_t6,N2533_t7,N2542_t0,
     N2542_t1,N2542_t2,N2542_t3,N2542_t4,N2542_t5,N2542_t6,N2542_t7,N2551_t0,N2551_t1,N2551_t2,
     N2551_t3,N2551_t4,N2551_t5,N2551_t6,N2551_t7,N2560_t0,N2560_t1,N2560_t2,N2560_t3,N2560_t4,
     N2560_t5,N2560_t6,N2560_t7,N2569_t0,N2569_t1,N2569_t2,N2569_t3,N2569_t4,N2569_t5,N2569_t6,
     N2569_t7,N2578_t0,N2578_t1,N2578_t2,N2578_t3,N2578_t4,N2578_t5,N2578_t6,N2578_t7,N2587_t0,
     N2587_t1,N2587_t2,N2587_t3,N2587_t4,N2587_t5,N2587_t6,N2587_t7,N2596_t0,N2596_t1,N2596_t2,
     N2596_t3,N2596_t4,N2596_t5,N2596_t6,N2596_t7,N2605_t0,N2605_t1,N2605_t2,N2605_t3,N2605_t4,
     N2605_t5,N2605_t6,N2605_t7,N2614_t0,N2614_t1,N2614_t2,N2614_t3,N2614_t4,N2614_t5,N2614_t6,
     N2614_t7,N2623_t0,N2623_t1,N2623_t2,N2623_t3,N2623_t4,N2623_t5,N2623_t6,N2623_t7,N2656_t0,
     N2656_t1,N2652_t0,N2652_t1,N2652_t2,N2659_t0,N2659_t1,N2670_t0,N2670_t1,N2666_t0,N2666_t1,
     N2666_t2,N2681_t0,N2681_t1,N2677_t0,N2677_t1,N2677_t2,N2692_t0,N2692_t1,N2692_t2,N2692_t3,
     N2688_t0,N2688_t1,N2688_t2,N2697_t0,N2697_t1,N2697_t2,N2697_t3,N2710_t0,N2710_t1,N2710_t2,
     N2710_t3,N2706_t0,N2706_t1,N2706_t2,N2723_t0,N2723_t1,N2723_t2,N2723_t3,N2719_t0,N2719_t1,
     N2719_t2,N1909_t0,N1909_t1,N2648_t0,N2648_t1,N2648_t2,N1913_t0,N1913_t1,N1913_t2,N2662_t0,
     N2662_t1,N2662_t2,N2673_t0,N2673_t1,N2673_t2,N2684_t0,N2684_t1,N2684_t2,N1922_t0,N1922_t1,
     N1922_t2,N2702_t0,N2702_t1,N2702_t2,N2715_t0,N2715_t1,N2715_t2,N143_t0,N143_t1,N143_t2,
     N143_t3,N143_t4,N143_t5,N137_t0,N137_t1,N137_t2,N137_t3,N137_t4,N132_t0,N132_t1,
     N132_t2,N132_t3,N128_t0,N128_t1,N128_t2,N125_t0,N125_t1,N311_t0,N311_t1,N311_t2,
     N311_t3,N311_t4,N317_t0,N317_t1,N317_t2,N317_t3,N322_t0,N322_t1,N322_t2,N326_t0,
     N326_t1,N2977_t0,N2977_t1,N2973_t0,N2973_t1,N2973_t2,N3112_t0,N3112_t1,N3115_t0,N3115_t1,
     N3119_t0,N3119_t1,N1875_t0,N1875_t1,N2073_t0,N2073_t1,N3128_t0,N3128_t1,N3131_t0,N3131_t1,
     N3135_t0,N3135_t1,N3138_t0,N3138_t1,N3142_t0,N3142_t1,N3145_t0,N3145_t1,N3149_t0,N3149_t1,
     N1895_t0,N1895_t1,N2093_t0,N2093_t1,N3158_t0,N3158_t1,N3161_t0,N3161_t1,N3165_t0,N3165_t1,
     N3168_t0,N3168_t1,N2967_t0,N2967_t1,N2970_t0,N2970_t1,N3172_t0,N3172_t1,N3175_t0,N3175_t1,
     N3178_t0,N3178_t1,N3181_t0,N3181_t1,N3184_t0,N3184_t1,N3187_t0,N3187_t1,N3478_t0,N3478_t1,
     N3481_t0,N3481_t1,N3487_t0,N3487_t1,N3484_t0,N3484_t1,N3472_t0,N3472_t1,N3475_t0,N3475_t1,
     N3407_t0,N3407_t1,N3410_t0,N3410_t1,N3415_t0,N3415_t1,N3415_t2,N3122_t0,N3122_t1,N3125_t0,
     N3125_t1,N3419_t0,N3419_t1,N3419_t2,N3423_t0,N3423_t1,N3426_t0,N3426_t1,N3431_t0,N3431_t1,
     N3434_t0,N3434_t1,N3439_t0,N3439_t1,N3442_t0,N3442_t1,N3447_t0,N3447_t1,N3447_t2,N3152_t0,
     N3152_t1,N3155_t0,N3155_t1,N3451_t0,N3451_t1,N3451_t2,N3455_t0,N3455_t1,N3458_t0,N3458_t1,
     N3463_t0,N3463_t1,N3466_t0,N3466_t1,N3493_t0,N3493_t1,N3496_t0,N3496_t1,N3499_t0,N3499_t1,
     N3502_t0,N3502_t1,N3505_t0,N3505_t1,N3511_t0,N3511_t1,N3517_t0,N3517_t1,N3520_t0,N3520_t1,
     N3523_t0,N3523_t1,N3514_t0,N3514_t1,N3384_t0,N3384_t1,N3490_t0,N3490_t1,N3508_t0,N3508_t1,
     N3700_t0,N3700_t1,N3697_t0,N3697_t1,N3645_t0,N3645_t1,N3648_t0,N3648_t1,N3664_t0,N3664_t1,
     N3667_t0,N3667_t1,N3654_t0,N3654_t1,N3658_t0,N3658_t1,N3673_t0,N3673_t1,N1926_t0,N1926_t1,
     N1926_t2,N3677_t0,N3677_t1,N3682_t0,N3682_t1,N3690_t0,N3690_t1,N3721_t0,N3721_t1,N3721_t2,
     N3721_t3,N3721_t4,N3734_t0,N3734_t1,N3734_t2,N3740_t0,N3740_t1,N3743_t0,N3743_t1,N3743_t2,
     N3743_t3,N3743_t4,N3756_t0,N3756_t1,N3756_t2,N3762_t0,N3762_t1,N3786_t0,N3786_t1,N3800_t0,
     N3800_t1,N3821_t0,N3821_t1,N3824_t0,N3824_t1,N3830_t0,N3830_t1,N3827_t0,N3827_t1,N3812_t0,
     N3812_t1,N3818_t0,N3818_t1,N3809_t0,N3809_t1,N3838_t0,N3838_t1,N3838_t2,N3838_t3,N3845_t0,
     N3845_t1,N3845_t2,N3845_t3,N3850_t0,N3850_t1,N3855_t0,N3855_t1,N3858_t0,N3858_t1,N3861_t0,
     N3861_t1,N3865_t0,N3865_t1,N3868_t0,N3868_t1,N3921_t0,N3921_t1,N3932_t0,N3932_t1,N3926_t0,
     N3926_t1,N3926_t2,N3953_t0,N3953_t1,N3959_t0,N3959_t1,N3965_t0,N3965_t1,N3971_t0,N3971_t1,
     N3977_t0,N3977_t1,N3983_t0,N3983_t1,N3956_t0,N3956_t1,N3962_t0,N3962_t1,N3980_t0,N3980_t1,
     N3974_t0,N3974_t1,N3950_t0,N3950_t1,N3937_t0,N3937_t1,N3968_t0,N3968_t1,N3940_t0,N3940_t1,
     N3996_t0,N3996_t1,N3992_t0,N3992_t1,N4062_t0,N4062_t1,N4070_t0,N4070_t1,N4059_t0,N4059_t1,
     N4067_t0,N4067_t1,N4091_t0,N4091_t1,N4094_t0,N4094_t1,N4094_t2,N4116_t0,N4116_t1,N4119_t0,
     N4119_t1,N4123_t0,N4123_t1,N4128_t0,N4128_t1,N4128_t2,N4128_t3,N4128_t4,N3917_t0,N3917_t1,
     N4139_t0,N4139_t1,N4142_t0,N4142_t1,N4167_t0,N4167_t1,N4167_t2,N4167_t3,N4167_t4,N4167_t5,
     N4035_t0,N4035_t1,N4174_t0,N4174_t1,N4174_t2,N4174_t3,N3815_t0,N3815_t1,N4186_t0,N4186_t1,
     N4182_t0,N4182_t1,N4197_t0,N4197_t1,N4213_t0,N4213_t1,N4213_t2,N4213_t3,N4203_t0,N4203_t1,
     N4203_t2,N4203_t3,N4203_t4,N4209_t0,N4209_t1,N4209_t2,N4223_t0,N4223_t1,N4223_t2,N4223_t3,
     N4218_t0,N4218_t1,N4218_t2,N4218_t3,N3913_t0,N3913_t1,N4247_t0,N4247_t1,N4242_t0,N4242_t1,
     N4287_t0,N4287_t1,N4287_t2,N4284_t0,N4284_t1,N4331_t0,N4331_t1,N4296_t0,N4296_t1,N4305_t0,
     N4305_t1,N4305_t2,N4305_t3,N4200_t0,N4200_t1,N4356_t0,N4356_t1,N4365_t0,N4365_t1,N4368_t0,
     N4368_t1,N4371_t0,N4371_t1,N4310_t0,N4310_t1,N4310_t2,N4353_t0,N4353_t1,N4359_t0,N4359_t1,
     N4362_t0,N4362_t1,N4319_t0,N4319_t1,N4398_t0,N4398_t1,N4413_t0,N4413_t1,N4435_t0,N4435_t1,
     N4421_t0,N4421_t1,N4427_t0,N4427_t1,N4416_t0,N4416_t1,N4430_t0,N4430_t1,N4387_t0,N4387_t1,
     N4390_t0,N4390_t1,N4443_t0,N4443_t1,N4493_t0,N4493_t1,N4465_t0,N4465_t1,N4468_t0,N4468_t1,
     N4479_t0,N4479_t1,N4458_t0,N4458_t1,N2758_t0,N2758_t1,N4498_t0,N4498_t1,N2761_t0,N2761_t1,
     N4531_t0,N4531_t1,N4534_t0,N4534_t1,N4537_t0,N4537_t1,N4540_t0,N4540_t1,N4503_t0,N4503_t1,
     N4569_t0,N4569_t1,N4576_t0,N4576_t1,N4581_t0,N4581_t1,N4584_t0,N4584_t1,N4559_t0,N4559_t1,
     N4549_t0,N4549_t1,N4564_t0,N4564_t1,N4564_t2,N4616_t0,N4616_t1,N4619_t0,N4619_t1,N4623_t0,
     N4623_t1,N4613_t0,N4613_t1,N4593_t0,N4593_t1,N4599_t0,N4599_t1,N4656_t0,N4656_t1,N4659_t0,
     N4659_t1,N4644_t0,N4644_t1,N4664_t0,N4664_t1,N4647_t0,N4647_t1,N4650_t0,N4650_t1,N4350_t0,
     N4350_t1,N4691_t0,N4691_t1,N4694_t0,N4694_t1,N4697_t0,N4697_t1,N4700_t0,N4700_t1,N4730_t0,
     N4730_t1,N4711_t0,N4711_t1,N4717_t0,N4717_t1,N4717_t2,N4722_t0,N4722_t1,N4722_t2,N4727_t0,
     N4727_t1,N4769_t0,N4769_t1,N4772_t0,N4772_t1,N4775_t0,N4775_t1,N4743_t0,N4743_t1,N4743_t2,
     N4757_t0,N4757_t1,N4757_t2,N4740_t0,N4740_t1,N4805_t0,N4805_t1,N4808_t0,N4808_t1,N4794_t0,
     N4794_t1,N4797_t0,N4797_t1,N4341_t0,N4341_t1,N4812_t0,N4812_t1,N4844_t0,N4844_t1,N4847_t0,
     N4847_t1,N4823_t0,N4823_t1,N4850_t0,N4850_t1,N4854_t0,N4854_t1,N4818_t0,N4818_t1,N4818_t2,
     N4880_t0,N4880_t1,N4889_t0,N4889_t1,N4876_t0,N4876_t1,N4876_t2,N4916_t0,N4916_t1,N2764_t0,
     N2764_t1,N2483_t0,N2483_t1,N4921_t0,N4921_t1,N4937_t0,N4937_t1,N4940_t0,N4940_t1,N4946_t0,
     N4946_t1,N4913_t0,N4913_t1,N4954_t0,N4954_t1,N4344_t0,N4344_t1,N4800_t0,N4800_t1,N4957_t0,
     N4957_t1,N4347_t0,N4347_t1,N4838_t0,N4838_t1,N4973_t0,N4973_t1,N4475_t0,N4475_t1,N4991_t0,
     N4991_t1,N4999_t0,N4999_t1,N4996_t0,N4996_t1,N4988_t0,N4988_t1,N5021_t0,N5021_t1,N4831_t0,
     N4831_t1,N5010_t0,N5010_t1,N4472_t0,N4472_t1,N4907_t0,N4907_t1,N5013_t0,N5013_t1,N4338_t0,
     N4338_t1,N5018_t0,N5018_t1,N4985_t0,N4985_t1,N5030_t0,N5030_t1,N4335_t0,N4335_t1,N5039_t0,
     N5039_t1,N5042_t0,N5042_t1,N5050_t0,N5050_t1,N5050_t2,N5050_t3,N5061_t0,N5061_t1,N5070_t0,
     N5070_t1,N5058_t0,N5058_t1,N1461_t0,N1461_t1,N5080_t0,N5080_t1,N5080_t2,N5080_t3,N5055_t0,
     N5055_t1,N5085_t0,N5085_t1,N5111_t0,N5111_t1,N5117_t0,N5117_t1,N5114_t0,N5114_t1,N5066_t0,
     N5066_t1,N5133_t0,N5133_t1,N5122_t0,N5122_t1,N5139_t0,N5139_t1,N5128_t0,N5128_t1,N5151_t0,
     N5151_t1,N5154_t0,N5154_t1,N5160_t0,N5160_t1,N5163_t0,N5163_t1,N5145_t0,N5145_t1,N5174_t0,
     N5174_t1,N5177_t0,N5177_t1,N5184_t0,N5184_t1,N5188_t0,N5188_t1,N5205_t0,N5205_t1,N5209_t0,
     N5209_t1,N5228_t0,N5228_t1,N5236_t0,N5236_t1,N5236_t2,N5254_t0,N5254_t1,N2307_t0,N2307_t1,
     N5250_t0,N5250_t1,N2310_t0,N2310_t1,N5269_t0,N5269_t1,N5266_t0,N5266_t1,N5258_t0,N5258_t1,
     N5279_t0,N5279_t1,N5292_t0,N5292_t1,N5289_t0,N5289_t1,N5306_t0,N5306_t1,N5303_t0,N5303_t1,
     N5298_t0,N5298_t1,N5309_t0,N5309_t1,N5324_t0,N5324_t1,N5327_t0,N5327_t1,N5332_t0,N5332_t1,
     N5335_t0,N5335_t1;
reg [1824:0] FEN;
fim PI_N124( .fault(fault), .net(N124), .FEN(FEN[0]), .op(N124_t) );
fim PI_N222( .fault(fault), .net(N222), .FEN(FEN[1]), .op(N222_t) );
fim PI_N329( .fault(fault), .net(N329), .FEN(FEN[2]), .op(N329_t) );
fim PI_N349( .fault(fault), .net(N349), .FEN(FEN[3]), .op(N349_t) );
fim FAN_N50_0 ( .fault(fault), .net(N50), .FEN(FEN[4]), .op(N50_t0) );
fim FAN_N50_1 ( .fault(fault), .net(N50), .FEN(FEN[5]), .op(N50_t1) );
fim FAN_N50_2 ( .fault(fault), .net(N50), .FEN(FEN[6]), .op(N50_t2) );
fim FAN_N50_3 ( .fault(fault), .net(N50), .FEN(FEN[7]), .op(N50_t3) );
fim FAN_N50_4 ( .fault(fault), .net(N50), .FEN(FEN[8]), .op(N50_t4) );
fim FAN_N50_5 ( .fault(fault), .net(N50), .FEN(FEN[9]), .op(N50_t5) );
fim FAN_N50_6 ( .fault(fault), .net(N50), .FEN(FEN[10]), .op(N50_t6) );
fim FAN_N58_0 ( .fault(fault), .net(N58), .FEN(FEN[11]), .op(N58_t0) );
fim FAN_N58_1 ( .fault(fault), .net(N58), .FEN(FEN[12]), .op(N58_t1) );
fim FAN_N58_2 ( .fault(fault), .net(N58), .FEN(FEN[13]), .op(N58_t2) );
fim FAN_N58_3 ( .fault(fault), .net(N58), .FEN(FEN[14]), .op(N58_t3) );
fim FAN_N58_4 ( .fault(fault), .net(N58), .FEN(FEN[15]), .op(N58_t4) );
fim FAN_N58_5 ( .fault(fault), .net(N58), .FEN(FEN[16]), .op(N58_t5) );
fim FAN_N58_6 ( .fault(fault), .net(N58), .FEN(FEN[17]), .op(N58_t6) );
fim FAN_N58_7 ( .fault(fault), .net(N58), .FEN(FEN[18]), .op(N58_t7) );
fim FAN_N58_8 ( .fault(fault), .net(N58), .FEN(FEN[19]), .op(N58_t8) );
fim FAN_N68_0 ( .fault(fault), .net(N68), .FEN(FEN[20]), .op(N68_t0) );
fim FAN_N68_1 ( .fault(fault), .net(N68), .FEN(FEN[21]), .op(N68_t1) );
fim FAN_N68_2 ( .fault(fault), .net(N68), .FEN(FEN[22]), .op(N68_t2) );
fim FAN_N68_3 ( .fault(fault), .net(N68), .FEN(FEN[23]), .op(N68_t3) );
fim FAN_N68_4 ( .fault(fault), .net(N68), .FEN(FEN[24]), .op(N68_t4) );
fim FAN_N68_5 ( .fault(fault), .net(N68), .FEN(FEN[25]), .op(N68_t5) );
fim FAN_N68_6 ( .fault(fault), .net(N68), .FEN(FEN[26]), .op(N68_t6) );
fim FAN_N68_7 ( .fault(fault), .net(N68), .FEN(FEN[27]), .op(N68_t7) );
fim FAN_N77_0 ( .fault(fault), .net(N77), .FEN(FEN[28]), .op(N77_t0) );
fim FAN_N77_1 ( .fault(fault), .net(N77), .FEN(FEN[29]), .op(N77_t1) );
fim FAN_N77_2 ( .fault(fault), .net(N77), .FEN(FEN[30]), .op(N77_t2) );
fim FAN_N77_3 ( .fault(fault), .net(N77), .FEN(FEN[31]), .op(N77_t3) );
fim FAN_N77_4 ( .fault(fault), .net(N77), .FEN(FEN[32]), .op(N77_t4) );
fim FAN_N77_5 ( .fault(fault), .net(N77), .FEN(FEN[33]), .op(N77_t5) );
fim FAN_N77_6 ( .fault(fault), .net(N77), .FEN(FEN[34]), .op(N77_t6) );
fim FAN_N77_7 ( .fault(fault), .net(N77), .FEN(FEN[35]), .op(N77_t7) );
fim FAN_N77_8 ( .fault(fault), .net(N77), .FEN(FEN[36]), .op(N77_t8) );
fim FAN_N87_0 ( .fault(fault), .net(N87), .FEN(FEN[37]), .op(N87_t0) );
fim FAN_N87_1 ( .fault(fault), .net(N87), .FEN(FEN[38]), .op(N87_t1) );
fim FAN_N87_2 ( .fault(fault), .net(N87), .FEN(FEN[39]), .op(N87_t2) );
fim FAN_N87_3 ( .fault(fault), .net(N87), .FEN(FEN[40]), .op(N87_t3) );
fim FAN_N87_4 ( .fault(fault), .net(N87), .FEN(FEN[41]), .op(N87_t4) );
fim FAN_N87_5 ( .fault(fault), .net(N87), .FEN(FEN[42]), .op(N87_t5) );
fim FAN_N87_6 ( .fault(fault), .net(N87), .FEN(FEN[43]), .op(N87_t6) );
fim FAN_N87_7 ( .fault(fault), .net(N87), .FEN(FEN[44]), .op(N87_t7) );
fim FAN_N87_8 ( .fault(fault), .net(N87), .FEN(FEN[45]), .op(N87_t8) );
fim FAN_N97_0 ( .fault(fault), .net(N97), .FEN(FEN[46]), .op(N97_t0) );
fim FAN_N97_1 ( .fault(fault), .net(N97), .FEN(FEN[47]), .op(N97_t1) );
fim FAN_N97_2 ( .fault(fault), .net(N97), .FEN(FEN[48]), .op(N97_t2) );
fim FAN_N97_3 ( .fault(fault), .net(N97), .FEN(FEN[49]), .op(N97_t3) );
fim FAN_N97_4 ( .fault(fault), .net(N97), .FEN(FEN[50]), .op(N97_t4) );
fim FAN_N97_5 ( .fault(fault), .net(N97), .FEN(FEN[51]), .op(N97_t5) );
fim FAN_N97_6 ( .fault(fault), .net(N97), .FEN(FEN[52]), .op(N97_t6) );
fim FAN_N97_7 ( .fault(fault), .net(N97), .FEN(FEN[53]), .op(N97_t7) );
fim FAN_N97_8 ( .fault(fault), .net(N97), .FEN(FEN[54]), .op(N97_t8) );
fim FAN_N107_0 ( .fault(fault), .net(N107), .FEN(FEN[55]), .op(N107_t0) );
fim FAN_N107_1 ( .fault(fault), .net(N107), .FEN(FEN[56]), .op(N107_t1) );
fim FAN_N107_2 ( .fault(fault), .net(N107), .FEN(FEN[57]), .op(N107_t2) );
fim FAN_N107_3 ( .fault(fault), .net(N107), .FEN(FEN[58]), .op(N107_t3) );
fim FAN_N107_4 ( .fault(fault), .net(N107), .FEN(FEN[59]), .op(N107_t4) );
fim FAN_N107_5 ( .fault(fault), .net(N107), .FEN(FEN[60]), .op(N107_t5) );
fim FAN_N107_6 ( .fault(fault), .net(N107), .FEN(FEN[61]), .op(N107_t6) );
fim FAN_N107_7 ( .fault(fault), .net(N107), .FEN(FEN[62]), .op(N107_t7) );
fim FAN_N116_0 ( .fault(fault), .net(N116), .FEN(FEN[63]), .op(N116_t0) );
fim FAN_N116_1 ( .fault(fault), .net(N116), .FEN(FEN[64]), .op(N116_t1) );
fim FAN_N116_2 ( .fault(fault), .net(N116), .FEN(FEN[65]), .op(N116_t2) );
fim FAN_N116_3 ( .fault(fault), .net(N116), .FEN(FEN[66]), .op(N116_t3) );
fim FAN_N116_4 ( .fault(fault), .net(N116), .FEN(FEN[67]), .op(N116_t4) );
fim FAN_N116_5 ( .fault(fault), .net(N116), .FEN(FEN[68]), .op(N116_t5) );
fim FAN_N116_6 ( .fault(fault), .net(N116), .FEN(FEN[69]), .op(N116_t6) );
fim FAN_N257_0 ( .fault(fault), .net(N257), .FEN(FEN[70]), .op(N257_t0) );
fim FAN_N257_1 ( .fault(fault), .net(N257), .FEN(FEN[71]), .op(N257_t1) );
fim FAN_N257_2 ( .fault(fault), .net(N257), .FEN(FEN[72]), .op(N257_t2) );
fim FAN_N257_3 ( .fault(fault), .net(N257), .FEN(FEN[73]), .op(N257_t3) );
fim FAN_N257_4 ( .fault(fault), .net(N257), .FEN(FEN[74]), .op(N257_t4) );
fim FAN_N257_5 ( .fault(fault), .net(N257), .FEN(FEN[75]), .op(N257_t5) );
fim FAN_N264_0 ( .fault(fault), .net(N264), .FEN(FEN[76]), .op(N264_t0) );
fim FAN_N264_1 ( .fault(fault), .net(N264), .FEN(FEN[77]), .op(N264_t1) );
fim FAN_N264_2 ( .fault(fault), .net(N264), .FEN(FEN[78]), .op(N264_t2) );
fim FAN_N264_3 ( .fault(fault), .net(N264), .FEN(FEN[79]), .op(N264_t3) );
fim FAN_N264_4 ( .fault(fault), .net(N264), .FEN(FEN[80]), .op(N264_t4) );
fim FAN_N1_0 ( .fault(fault), .net(N1), .FEN(FEN[81]), .op(N1_t0) );
fim FAN_N1_1 ( .fault(fault), .net(N1), .FEN(FEN[82]), .op(N1_t1) );
fim FAN_N1_2 ( .fault(fault), .net(N1), .FEN(FEN[83]), .op(N1_t2) );
fim FAN_N1_3 ( .fault(fault), .net(N1), .FEN(FEN[84]), .op(N1_t3) );
fim FAN_N1_4 ( .fault(fault), .net(N1), .FEN(FEN[85]), .op(N1_t4) );
fim FAN_N1_5 ( .fault(fault), .net(N1), .FEN(FEN[86]), .op(N1_t5) );
fim FAN_N1_6 ( .fault(fault), .net(N1), .FEN(FEN[87]), .op(N1_t6) );
fim FAN_N1_7 ( .fault(fault), .net(N1), .FEN(FEN[88]), .op(N1_t7) );
fim FAN_N1_8 ( .fault(fault), .net(N1), .FEN(FEN[89]), .op(N1_t8) );
fim FAN_N1_9 ( .fault(fault), .net(N1), .FEN(FEN[90]), .op(N1_t9) );
fim FAN_N1_10 ( .fault(fault), .net(N1), .FEN(FEN[91]), .op(N1_t10) );
fim FAN_N13_0 ( .fault(fault), .net(N13), .FEN(FEN[92]), .op(N13_t0) );
fim FAN_N13_1 ( .fault(fault), .net(N13), .FEN(FEN[93]), .op(N13_t1) );
fim FAN_N13_2 ( .fault(fault), .net(N13), .FEN(FEN[94]), .op(N13_t2) );
fim FAN_N13_3 ( .fault(fault), .net(N13), .FEN(FEN[95]), .op(N13_t3) );
fim FAN_N13_4 ( .fault(fault), .net(N13), .FEN(FEN[96]), .op(N13_t4) );
fim FAN_N13_5 ( .fault(fault), .net(N13), .FEN(FEN[97]), .op(N13_t5) );
fim FAN_N20_0 ( .fault(fault), .net(N20), .FEN(FEN[98]), .op(N20_t0) );
fim FAN_N20_1 ( .fault(fault), .net(N20), .FEN(FEN[99]), .op(N20_t1) );
fim FAN_N20_2 ( .fault(fault), .net(N20), .FEN(FEN[100]), .op(N20_t2) );
fim FAN_N20_3 ( .fault(fault), .net(N20), .FEN(FEN[101]), .op(N20_t3) );
fim FAN_N20_4 ( .fault(fault), .net(N20), .FEN(FEN[102]), .op(N20_t4) );
fim FAN_N20_5 ( .fault(fault), .net(N20), .FEN(FEN[103]), .op(N20_t5) );
fim FAN_N20_6 ( .fault(fault), .net(N20), .FEN(FEN[104]), .op(N20_t6) );
fim FAN_N20_7 ( .fault(fault), .net(N20), .FEN(FEN[105]), .op(N20_t7) );
fim FAN_N20_8 ( .fault(fault), .net(N20), .FEN(FEN[106]), .op(N20_t8) );
fim FAN_N20_9 ( .fault(fault), .net(N20), .FEN(FEN[107]), .op(N20_t9) );
fim FAN_N20_10 ( .fault(fault), .net(N20), .FEN(FEN[108]), .op(N20_t10) );
fim FAN_N20_11 ( .fault(fault), .net(N20), .FEN(FEN[109]), .op(N20_t11) );
fim FAN_N33_0 ( .fault(fault), .net(N33), .FEN(FEN[110]), .op(N33_t0) );
fim FAN_N33_1 ( .fault(fault), .net(N33), .FEN(FEN[111]), .op(N33_t1) );
fim FAN_N33_2 ( .fault(fault), .net(N33), .FEN(FEN[112]), .op(N33_t2) );
fim FAN_N33_3 ( .fault(fault), .net(N33), .FEN(FEN[113]), .op(N33_t3) );
fim FAN_N33_4 ( .fault(fault), .net(N33), .FEN(FEN[114]), .op(N33_t4) );
fim FAN_N33_5 ( .fault(fault), .net(N33), .FEN(FEN[115]), .op(N33_t5) );
fim FAN_N33_6 ( .fault(fault), .net(N33), .FEN(FEN[116]), .op(N33_t6) );
fim FAN_N41_0 ( .fault(fault), .net(N41), .FEN(FEN[117]), .op(N41_t0) );
fim FAN_N41_1 ( .fault(fault), .net(N41), .FEN(FEN[118]), .op(N41_t1) );
fim FAN_N41_2 ( .fault(fault), .net(N41), .FEN(FEN[119]), .op(N41_t2) );
fim FAN_N45_0 ( .fault(fault), .net(N45), .FEN(FEN[120]), .op(N45_t0) );
fim FAN_N45_1 ( .fault(fault), .net(N45), .FEN(FEN[121]), .op(N45_t1) );
fim FAN_N45_2 ( .fault(fault), .net(N45), .FEN(FEN[122]), .op(N45_t2) );
fim FAN_N45_3 ( .fault(fault), .net(N45), .FEN(FEN[123]), .op(N45_t3) );
fim FAN_N190_0 ( .fault(fault), .net(N190), .FEN(FEN[124]), .op(N190_t0) );
fim FAN_N190_1 ( .fault(fault), .net(N190), .FEN(FEN[125]), .op(N190_t1) );
fim FAN_N190_2 ( .fault(fault), .net(N190), .FEN(FEN[126]), .op(N190_t2) );
fim FAN_N190_3 ( .fault(fault), .net(N190), .FEN(FEN[127]), .op(N190_t3) );
fim FAN_N190_4 ( .fault(fault), .net(N190), .FEN(FEN[128]), .op(N190_t4) );
fim FAN_N190_5 ( .fault(fault), .net(N190), .FEN(FEN[129]), .op(N190_t5) );
fim FAN_N190_6 ( .fault(fault), .net(N190), .FEN(FEN[130]), .op(N190_t6) );
fim FAN_N190_7 ( .fault(fault), .net(N190), .FEN(FEN[131]), .op(N190_t7) );
fim FAN_N190_8 ( .fault(fault), .net(N190), .FEN(FEN[132]), .op(N190_t8) );
fim FAN_N200_0 ( .fault(fault), .net(N200), .FEN(FEN[133]), .op(N200_t0) );
fim FAN_N200_1 ( .fault(fault), .net(N200), .FEN(FEN[134]), .op(N200_t1) );
fim FAN_N200_2 ( .fault(fault), .net(N200), .FEN(FEN[135]), .op(N200_t2) );
fim FAN_N200_3 ( .fault(fault), .net(N200), .FEN(FEN[136]), .op(N200_t3) );
fim FAN_N200_4 ( .fault(fault), .net(N200), .FEN(FEN[137]), .op(N200_t4) );
fim FAN_N200_5 ( .fault(fault), .net(N200), .FEN(FEN[138]), .op(N200_t5) );
fim FAN_N200_6 ( .fault(fault), .net(N200), .FEN(FEN[139]), .op(N200_t6) );
fim FAN_N200_7 ( .fault(fault), .net(N200), .FEN(FEN[140]), .op(N200_t7) );
fim FAN_N200_8 ( .fault(fault), .net(N200), .FEN(FEN[141]), .op(N200_t8) );
fim FAN_N200_9 ( .fault(fault), .net(N200), .FEN(FEN[142]), .op(N200_t9) );
fim FAN_N200_10 ( .fault(fault), .net(N200), .FEN(FEN[143]), .op(N200_t10) );
fim FAN_N200_11 ( .fault(fault), .net(N200), .FEN(FEN[144]), .op(N200_t11) );
fim FAN_N179_0 ( .fault(fault), .net(N179), .FEN(FEN[145]), .op(N179_t0) );
fim FAN_N179_1 ( .fault(fault), .net(N179), .FEN(FEN[146]), .op(N179_t1) );
fim FAN_N179_2 ( .fault(fault), .net(N179), .FEN(FEN[147]), .op(N179_t2) );
fim FAN_N179_3 ( .fault(fault), .net(N179), .FEN(FEN[148]), .op(N179_t3) );
fim FAN_N179_4 ( .fault(fault), .net(N179), .FEN(FEN[149]), .op(N179_t4) );
fim FAN_N179_5 ( .fault(fault), .net(N179), .FEN(FEN[150]), .op(N179_t5) );
fim FAN_N179_6 ( .fault(fault), .net(N179), .FEN(FEN[151]), .op(N179_t6) );
fim FAN_N179_7 ( .fault(fault), .net(N179), .FEN(FEN[152]), .op(N179_t7) );
fim FAN_N179_8 ( .fault(fault), .net(N179), .FEN(FEN[153]), .op(N179_t8) );
fim FAN_N179_9 ( .fault(fault), .net(N179), .FEN(FEN[154]), .op(N179_t9) );
fim FAN_N213_0 ( .fault(fault), .net(N213), .FEN(FEN[155]), .op(N213_t0) );
fim FAN_N213_1 ( .fault(fault), .net(N213), .FEN(FEN[156]), .op(N213_t1) );
fim FAN_N213_2 ( .fault(fault), .net(N213), .FEN(FEN[157]), .op(N213_t2) );
fim FAN_N213_3 ( .fault(fault), .net(N213), .FEN(FEN[158]), .op(N213_t3) );
fim FAN_N213_4 ( .fault(fault), .net(N213), .FEN(FEN[159]), .op(N213_t4) );
fim FAN_N213_5 ( .fault(fault), .net(N213), .FEN(FEN[160]), .op(N213_t5) );
fim FAN_N213_6 ( .fault(fault), .net(N213), .FEN(FEN[161]), .op(N213_t6) );
fim FAN_N213_7 ( .fault(fault), .net(N213), .FEN(FEN[162]), .op(N213_t7) );
fim FAN_N343_0 ( .fault(fault), .net(N343), .FEN(FEN[163]), .op(N343_t0) );
fim FAN_N343_1 ( .fault(fault), .net(N343), .FEN(FEN[164]), .op(N343_t1) );
fim FAN_N343_2 ( .fault(fault), .net(N343), .FEN(FEN[165]), .op(N343_t2) );
fim FAN_N343_3 ( .fault(fault), .net(N343), .FEN(FEN[166]), .op(N343_t3) );
fim FAN_N343_4 ( .fault(fault), .net(N343), .FEN(FEN[167]), .op(N343_t4) );
fim FAN_N226_0 ( .fault(fault), .net(N226), .FEN(FEN[168]), .op(N226_t0) );
fim FAN_N226_1 ( .fault(fault), .net(N226), .FEN(FEN[169]), .op(N226_t1) );
fim FAN_N226_2 ( .fault(fault), .net(N226), .FEN(FEN[170]), .op(N226_t2) );
fim FAN_N226_3 ( .fault(fault), .net(N226), .FEN(FEN[171]), .op(N226_t3) );
fim FAN_N226_4 ( .fault(fault), .net(N226), .FEN(FEN[172]), .op(N226_t4) );
fim FAN_N232_0 ( .fault(fault), .net(N232), .FEN(FEN[173]), .op(N232_t0) );
fim FAN_N232_1 ( .fault(fault), .net(N232), .FEN(FEN[174]), .op(N232_t1) );
fim FAN_N232_2 ( .fault(fault), .net(N232), .FEN(FEN[175]), .op(N232_t2) );
fim FAN_N232_3 ( .fault(fault), .net(N232), .FEN(FEN[176]), .op(N232_t3) );
fim FAN_N232_4 ( .fault(fault), .net(N232), .FEN(FEN[177]), .op(N232_t4) );
fim FAN_N238_0 ( .fault(fault), .net(N238), .FEN(FEN[178]), .op(N238_t0) );
fim FAN_N238_1 ( .fault(fault), .net(N238), .FEN(FEN[179]), .op(N238_t1) );
fim FAN_N238_2 ( .fault(fault), .net(N238), .FEN(FEN[180]), .op(N238_t2) );
fim FAN_N238_3 ( .fault(fault), .net(N238), .FEN(FEN[181]), .op(N238_t3) );
fim FAN_N238_4 ( .fault(fault), .net(N238), .FEN(FEN[182]), .op(N238_t4) );
fim FAN_N244_0 ( .fault(fault), .net(N244), .FEN(FEN[183]), .op(N244_t0) );
fim FAN_N244_1 ( .fault(fault), .net(N244), .FEN(FEN[184]), .op(N244_t1) );
fim FAN_N244_2 ( .fault(fault), .net(N244), .FEN(FEN[185]), .op(N244_t2) );
fim FAN_N244_3 ( .fault(fault), .net(N244), .FEN(FEN[186]), .op(N244_t3) );
fim FAN_N244_4 ( .fault(fault), .net(N244), .FEN(FEN[187]), .op(N244_t4) );
fim FAN_N250_0 ( .fault(fault), .net(N250), .FEN(FEN[188]), .op(N250_t0) );
fim FAN_N250_1 ( .fault(fault), .net(N250), .FEN(FEN[189]), .op(N250_t1) );
fim FAN_N250_2 ( .fault(fault), .net(N250), .FEN(FEN[190]), .op(N250_t2) );
fim FAN_N250_3 ( .fault(fault), .net(N250), .FEN(FEN[191]), .op(N250_t3) );
fim FAN_N250_4 ( .fault(fault), .net(N250), .FEN(FEN[192]), .op(N250_t4) );
fim FAN_N250_5 ( .fault(fault), .net(N250), .FEN(FEN[193]), .op(N250_t5) );
fim FAN_N270_0 ( .fault(fault), .net(N270), .FEN(FEN[194]), .op(N270_t0) );
fim FAN_N270_1 ( .fault(fault), .net(N270), .FEN(FEN[195]), .op(N270_t1) );
fim FAN_N270_2 ( .fault(fault), .net(N270), .FEN(FEN[196]), .op(N270_t2) );
fim FAN_N330_0 ( .fault(fault), .net(N330), .FEN(FEN[197]), .op(N330_t0) );
fim FAN_N330_1 ( .fault(fault), .net(N330), .FEN(FEN[198]), .op(N330_t1) );
fim FAN_N330_2 ( .fault(fault), .net(N330), .FEN(FEN[199]), .op(N330_t2) );
fim FAN_N330_3 ( .fault(fault), .net(N330), .FEN(FEN[200]), .op(N330_t3) );
fim FAN_N330_4 ( .fault(fault), .net(N330), .FEN(FEN[201]), .op(N330_t4) );
fim FAN_N330_5 ( .fault(fault), .net(N330), .FEN(FEN[202]), .op(N330_t5) );
fim FAN_N330_6 ( .fault(fault), .net(N330), .FEN(FEN[203]), .op(N330_t6) );
fim FAN_N330_7 ( .fault(fault), .net(N330), .FEN(FEN[204]), .op(N330_t7) );
fim FAN_N330_8 ( .fault(fault), .net(N330), .FEN(FEN[205]), .op(N330_t8) );
fim FAN_N330_9 ( .fault(fault), .net(N330), .FEN(FEN[206]), .op(N330_t9) );
fim FAN_N330_10 ( .fault(fault), .net(N330), .FEN(FEN[207]), .op(N330_t10) );
fim FAN_N330_11 ( .fault(fault), .net(N330), .FEN(FEN[208]), .op(N330_t11) );
fim FAN_N169_0 ( .fault(fault), .net(N169), .FEN(FEN[209]), .op(N169_t0) );
fim FAN_N169_1 ( .fault(fault), .net(N169), .FEN(FEN[210]), .op(N169_t1) );
fim FAN_N169_2 ( .fault(fault), .net(N169), .FEN(FEN[211]), .op(N169_t2) );
fim FAN_N169_3 ( .fault(fault), .net(N169), .FEN(FEN[212]), .op(N169_t3) );
fim FAN_N169_4 ( .fault(fault), .net(N169), .FEN(FEN[213]), .op(N169_t4) );
fim FAN_N169_5 ( .fault(fault), .net(N169), .FEN(FEN[214]), .op(N169_t5) );
fim FAN_N169_6 ( .fault(fault), .net(N169), .FEN(FEN[215]), .op(N169_t6) );
fim FAN_N169_7 ( .fault(fault), .net(N169), .FEN(FEN[216]), .op(N169_t7) );
fim FAN_N169_8 ( .fault(fault), .net(N169), .FEN(FEN[217]), .op(N169_t8) );
fim FAN_N842_0 ( .fault(fault), .net(N842), .FEN(FEN[218]), .op(N842_t0) );
fim FAN_N842_1 ( .fault(fault), .net(N842), .FEN(FEN[219]), .op(N842_t1) );
fim FAN_N848_0 ( .fault(fault), .net(N848), .FEN(FEN[220]), .op(N848_t0) );
fim FAN_N848_1 ( .fault(fault), .net(N848), .FEN(FEN[221]), .op(N848_t1) );
fim FAN_N854_0 ( .fault(fault), .net(N854), .FEN(FEN[222]), .op(N854_t0) );
fim FAN_N854_1 ( .fault(fault), .net(N854), .FEN(FEN[223]), .op(N854_t1) );
fim FAN_N854_2 ( .fault(fault), .net(N854), .FEN(FEN[224]), .op(N854_t2) );
fim FAN_N655_0 ( .fault(fault), .net(N655), .FEN(FEN[225]), .op(N655_t0) );
fim FAN_N655_1 ( .fault(fault), .net(N655), .FEN(FEN[226]), .op(N655_t1) );
fim FAN_N655_2 ( .fault(fault), .net(N655), .FEN(FEN[227]), .op(N655_t2) );
fim FAN_N655_3 ( .fault(fault), .net(N655), .FEN(FEN[228]), .op(N655_t3) );
fim FAN_N655_4 ( .fault(fault), .net(N655), .FEN(FEN[229]), .op(N655_t4) );
fim FAN_N655_5 ( .fault(fault), .net(N655), .FEN(FEN[230]), .op(N655_t5) );
fim FAN_N655_6 ( .fault(fault), .net(N655), .FEN(FEN[231]), .op(N655_t6) );
fim FAN_N655_7 ( .fault(fault), .net(N655), .FEN(FEN[232]), .op(N655_t7) );
fim FAN_N655_8 ( .fault(fault), .net(N655), .FEN(FEN[233]), .op(N655_t8) );
fim FAN_N670_0 ( .fault(fault), .net(N670), .FEN(FEN[234]), .op(N670_t0) );
fim FAN_N670_1 ( .fault(fault), .net(N670), .FEN(FEN[235]), .op(N670_t1) );
fim FAN_N670_2 ( .fault(fault), .net(N670), .FEN(FEN[236]), .op(N670_t2) );
fim FAN_N670_3 ( .fault(fault), .net(N670), .FEN(FEN[237]), .op(N670_t3) );
fim FAN_N670_4 ( .fault(fault), .net(N670), .FEN(FEN[238]), .op(N670_t4) );
fim FAN_N670_5 ( .fault(fault), .net(N670), .FEN(FEN[239]), .op(N670_t5) );
fim FAN_N670_6 ( .fault(fault), .net(N670), .FEN(FEN[240]), .op(N670_t6) );
fim FAN_N670_7 ( .fault(fault), .net(N670), .FEN(FEN[241]), .op(N670_t7) );
fim FAN_N690_0 ( .fault(fault), .net(N690), .FEN(FEN[242]), .op(N690_t0) );
fim FAN_N690_1 ( .fault(fault), .net(N690), .FEN(FEN[243]), .op(N690_t1) );
fim FAN_N690_2 ( .fault(fault), .net(N690), .FEN(FEN[244]), .op(N690_t2) );
fim FAN_N690_3 ( .fault(fault), .net(N690), .FEN(FEN[245]), .op(N690_t3) );
fim FAN_N690_4 ( .fault(fault), .net(N690), .FEN(FEN[246]), .op(N690_t4) );
fim FAN_N690_5 ( .fault(fault), .net(N690), .FEN(FEN[247]), .op(N690_t5) );
fim FAN_N690_6 ( .fault(fault), .net(N690), .FEN(FEN[248]), .op(N690_t6) );
fim FAN_N690_7 ( .fault(fault), .net(N690), .FEN(FEN[249]), .op(N690_t7) );
fim FAN_N706_0 ( .fault(fault), .net(N706), .FEN(FEN[250]), .op(N706_t0) );
fim FAN_N706_1 ( .fault(fault), .net(N706), .FEN(FEN[251]), .op(N706_t1) );
fim FAN_N706_2 ( .fault(fault), .net(N706), .FEN(FEN[252]), .op(N706_t2) );
fim FAN_N706_3 ( .fault(fault), .net(N706), .FEN(FEN[253]), .op(N706_t3) );
fim FAN_N706_4 ( .fault(fault), .net(N706), .FEN(FEN[254]), .op(N706_t4) );
fim FAN_N706_5 ( .fault(fault), .net(N706), .FEN(FEN[255]), .op(N706_t5) );
fim FAN_N706_6 ( .fault(fault), .net(N706), .FEN(FEN[256]), .op(N706_t6) );
fim FAN_N706_7 ( .fault(fault), .net(N706), .FEN(FEN[257]), .op(N706_t7) );
fim FAN_N715_0 ( .fault(fault), .net(N715), .FEN(FEN[258]), .op(N715_t0) );
fim FAN_N715_1 ( .fault(fault), .net(N715), .FEN(FEN[259]), .op(N715_t1) );
fim FAN_N715_2 ( .fault(fault), .net(N715), .FEN(FEN[260]), .op(N715_t2) );
fim FAN_N715_3 ( .fault(fault), .net(N715), .FEN(FEN[261]), .op(N715_t3) );
fim FAN_N715_4 ( .fault(fault), .net(N715), .FEN(FEN[262]), .op(N715_t4) );
fim FAN_N715_5 ( .fault(fault), .net(N715), .FEN(FEN[263]), .op(N715_t5) );
fim FAN_N715_6 ( .fault(fault), .net(N715), .FEN(FEN[264]), .op(N715_t6) );
fim FAN_N715_7 ( .fault(fault), .net(N715), .FEN(FEN[265]), .op(N715_t7) );
fim FAN_N727_0 ( .fault(fault), .net(N727), .FEN(FEN[266]), .op(N727_t0) );
fim FAN_N727_1 ( .fault(fault), .net(N727), .FEN(FEN[267]), .op(N727_t1) );
fim FAN_N727_2 ( .fault(fault), .net(N727), .FEN(FEN[268]), .op(N727_t2) );
fim FAN_N727_3 ( .fault(fault), .net(N727), .FEN(FEN[269]), .op(N727_t3) );
fim FAN_N727_4 ( .fault(fault), .net(N727), .FEN(FEN[270]), .op(N727_t4) );
fim FAN_N727_5 ( .fault(fault), .net(N727), .FEN(FEN[271]), .op(N727_t5) );
fim FAN_N727_6 ( .fault(fault), .net(N727), .FEN(FEN[272]), .op(N727_t6) );
fim FAN_N727_7 ( .fault(fault), .net(N727), .FEN(FEN[273]), .op(N727_t7) );
fim FAN_N740_0 ( .fault(fault), .net(N740), .FEN(FEN[274]), .op(N740_t0) );
fim FAN_N740_1 ( .fault(fault), .net(N740), .FEN(FEN[275]), .op(N740_t1) );
fim FAN_N740_2 ( .fault(fault), .net(N740), .FEN(FEN[276]), .op(N740_t2) );
fim FAN_N740_3 ( .fault(fault), .net(N740), .FEN(FEN[277]), .op(N740_t3) );
fim FAN_N740_4 ( .fault(fault), .net(N740), .FEN(FEN[278]), .op(N740_t4) );
fim FAN_N740_5 ( .fault(fault), .net(N740), .FEN(FEN[279]), .op(N740_t5) );
fim FAN_N740_6 ( .fault(fault), .net(N740), .FEN(FEN[280]), .op(N740_t6) );
fim FAN_N740_7 ( .fault(fault), .net(N740), .FEN(FEN[281]), .op(N740_t7) );
fim FAN_N753_0 ( .fault(fault), .net(N753), .FEN(FEN[282]), .op(N753_t0) );
fim FAN_N753_1 ( .fault(fault), .net(N753), .FEN(FEN[283]), .op(N753_t1) );
fim FAN_N753_2 ( .fault(fault), .net(N753), .FEN(FEN[284]), .op(N753_t2) );
fim FAN_N753_3 ( .fault(fault), .net(N753), .FEN(FEN[285]), .op(N753_t3) );
fim FAN_N753_4 ( .fault(fault), .net(N753), .FEN(FEN[286]), .op(N753_t4) );
fim FAN_N753_5 ( .fault(fault), .net(N753), .FEN(FEN[287]), .op(N753_t5) );
fim FAN_N753_6 ( .fault(fault), .net(N753), .FEN(FEN[288]), .op(N753_t6) );
fim FAN_N753_7 ( .fault(fault), .net(N753), .FEN(FEN[289]), .op(N753_t7) );
fim FAN_N753_8 ( .fault(fault), .net(N753), .FEN(FEN[290]), .op(N753_t8) );
fim FAN_N926_0 ( .fault(fault), .net(N926), .FEN(FEN[291]), .op(N926_t0) );
fim FAN_N926_1 ( .fault(fault), .net(N926), .FEN(FEN[292]), .op(N926_t1) );
fim FAN_N929_0 ( .fault(fault), .net(N929), .FEN(FEN[293]), .op(N929_t0) );
fim FAN_N929_1 ( .fault(fault), .net(N929), .FEN(FEN[294]), .op(N929_t1) );
fim FAN_N932_0 ( .fault(fault), .net(N932), .FEN(FEN[295]), .op(N932_t0) );
fim FAN_N932_1 ( .fault(fault), .net(N932), .FEN(FEN[296]), .op(N932_t1) );
fim FAN_N935_0 ( .fault(fault), .net(N935), .FEN(FEN[297]), .op(N935_t0) );
fim FAN_N935_1 ( .fault(fault), .net(N935), .FEN(FEN[298]), .op(N935_t1) );
fim FAN_N679_0 ( .fault(fault), .net(N679), .FEN(FEN[299]), .op(N679_t0) );
fim FAN_N679_1 ( .fault(fault), .net(N679), .FEN(FEN[300]), .op(N679_t1) );
fim FAN_N679_2 ( .fault(fault), .net(N679), .FEN(FEN[301]), .op(N679_t2) );
fim FAN_N686_0 ( .fault(fault), .net(N686), .FEN(FEN[302]), .op(N686_t0) );
fim FAN_N686_1 ( .fault(fault), .net(N686), .FEN(FEN[303]), .op(N686_t1) );
fim FAN_N686_2 ( .fault(fault), .net(N686), .FEN(FEN[304]), .op(N686_t2) );
fim FAN_N736_0 ( .fault(fault), .net(N736), .FEN(FEN[305]), .op(N736_t0) );
fim FAN_N736_1 ( .fault(fault), .net(N736), .FEN(FEN[306]), .op(N736_t1) );
fim FAN_N736_2 ( .fault(fault), .net(N736), .FEN(FEN[307]), .op(N736_t2) );
fim FAN_N749_0 ( .fault(fault), .net(N749), .FEN(FEN[308]), .op(N749_t0) );
fim FAN_N749_1 ( .fault(fault), .net(N749), .FEN(FEN[309]), .op(N749_t1) );
fim FAN_N749_2 ( .fault(fault), .net(N749), .FEN(FEN[310]), .op(N749_t2) );
fim FAN_N683_0 ( .fault(fault), .net(N683), .FEN(FEN[311]), .op(N683_t0) );
fim FAN_N683_1 ( .fault(fault), .net(N683), .FEN(FEN[312]), .op(N683_t1) );
fim FAN_N699_0 ( .fault(fault), .net(N699), .FEN(FEN[313]), .op(N699_t0) );
fim FAN_N699_1 ( .fault(fault), .net(N699), .FEN(FEN[314]), .op(N699_t1) );
fim FAN_N665_0 ( .fault(fault), .net(N665), .FEN(FEN[315]), .op(N665_t0) );
fim FAN_N665_1 ( .fault(fault), .net(N665), .FEN(FEN[316]), .op(N665_t1) );
fim FAN_N665_2 ( .fault(fault), .net(N665), .FEN(FEN[317]), .op(N665_t2) );
fim FAN_N665_3 ( .fault(fault), .net(N665), .FEN(FEN[318]), .op(N665_t3) );
fim FAN_N953_0 ( .fault(fault), .net(N953), .FEN(FEN[319]), .op(N953_t0) );
fim FAN_N953_1 ( .fault(fault), .net(N953), .FEN(FEN[320]), .op(N953_t1) );
fim FAN_N959_0 ( .fault(fault), .net(N959), .FEN(FEN[321]), .op(N959_t0) );
fim FAN_N959_1 ( .fault(fault), .net(N959), .FEN(FEN[322]), .op(N959_t1) );
fim FAN_N839_0 ( .fault(fault), .net(N839), .FEN(FEN[323]), .op(N839_t0) );
fim FAN_N839_1 ( .fault(fault), .net(N839), .FEN(FEN[324]), .op(N839_t1) );
fim FAN_N782_0 ( .fault(fault), .net(N782), .FEN(FEN[325]), .op(N782_t0) );
fim FAN_N782_1 ( .fault(fault), .net(N782), .FEN(FEN[326]), .op(N782_t1) );
fim FAN_N782_2 ( .fault(fault), .net(N782), .FEN(FEN[327]), .op(N782_t2) );
fim FAN_N825_0 ( .fault(fault), .net(N825), .FEN(FEN[328]), .op(N825_t0) );
fim FAN_N825_1 ( .fault(fault), .net(N825), .FEN(FEN[329]), .op(N825_t1) );
fim FAN_N825_2 ( .fault(fault), .net(N825), .FEN(FEN[330]), .op(N825_t2) );
fim FAN_N832_0 ( .fault(fault), .net(N832), .FEN(FEN[331]), .op(N832_t0) );
fim FAN_N832_1 ( .fault(fault), .net(N832), .FEN(FEN[332]), .op(N832_t1) );
fim FAN_N779_0 ( .fault(fault), .net(N779), .FEN(FEN[333]), .op(N779_t0) );
fim FAN_N779_1 ( .fault(fault), .net(N779), .FEN(FEN[334]), .op(N779_t1) );
fim FAN_N836_0 ( .fault(fault), .net(N836), .FEN(FEN[335]), .op(N836_t0) );
fim FAN_N836_1 ( .fault(fault), .net(N836), .FEN(FEN[336]), .op(N836_t1) );
fim FAN_N769_0 ( .fault(fault), .net(N769), .FEN(FEN[337]), .op(N769_t0) );
fim FAN_N769_1 ( .fault(fault), .net(N769), .FEN(FEN[338]), .op(N769_t1) );
fim FAN_N772_0 ( .fault(fault), .net(N772), .FEN(FEN[339]), .op(N772_t0) );
fim FAN_N772_1 ( .fault(fault), .net(N772), .FEN(FEN[340]), .op(N772_t1) );
fim FAN_N772_2 ( .fault(fault), .net(N772), .FEN(FEN[341]), .op(N772_t2) );
fim FAN_N772_3 ( .fault(fault), .net(N772), .FEN(FEN[342]), .op(N772_t3) );
fim FAN_N772_4 ( .fault(fault), .net(N772), .FEN(FEN[343]), .op(N772_t4) );
fim FAN_N772_5 ( .fault(fault), .net(N772), .FEN(FEN[344]), .op(N772_t5) );
fim FAN_N786_0 ( .fault(fault), .net(N786), .FEN(FEN[345]), .op(N786_t0) );
fim FAN_N786_1 ( .fault(fault), .net(N786), .FEN(FEN[346]), .op(N786_t1) );
fim FAN_N786_2 ( .fault(fault), .net(N786), .FEN(FEN[347]), .op(N786_t2) );
fim FAN_N786_3 ( .fault(fault), .net(N786), .FEN(FEN[348]), .op(N786_t3) );
fim FAN_N786_4 ( .fault(fault), .net(N786), .FEN(FEN[349]), .op(N786_t4) );
fim FAN_N786_5 ( .fault(fault), .net(N786), .FEN(FEN[350]), .op(N786_t5) );
fim FAN_N798_0 ( .fault(fault), .net(N798), .FEN(FEN[351]), .op(N798_t0) );
fim FAN_N798_1 ( .fault(fault), .net(N798), .FEN(FEN[352]), .op(N798_t1) );
fim FAN_N798_2 ( .fault(fault), .net(N798), .FEN(FEN[353]), .op(N798_t2) );
fim FAN_N798_3 ( .fault(fault), .net(N798), .FEN(FEN[354]), .op(N798_t3) );
fim FAN_N874_0 ( .fault(fault), .net(N874), .FEN(FEN[355]), .op(N874_t0) );
fim FAN_N874_1 ( .fault(fault), .net(N874), .FEN(FEN[356]), .op(N874_t1) );
fim FAN_N794_0 ( .fault(fault), .net(N794), .FEN(FEN[357]), .op(N794_t0) );
fim FAN_N794_1 ( .fault(fault), .net(N794), .FEN(FEN[358]), .op(N794_t1) );
fim FAN_N794_2 ( .fault(fault), .net(N794), .FEN(FEN[359]), .op(N794_t2) );
fim FAN_N956_0 ( .fault(fault), .net(N956), .FEN(FEN[360]), .op(N956_t0) );
fim FAN_N956_1 ( .fault(fault), .net(N956), .FEN(FEN[361]), .op(N956_t1) );
fim FAN_N861_0 ( .fault(fault), .net(N861), .FEN(FEN[362]), .op(N861_t0) );
fim FAN_N861_1 ( .fault(fault), .net(N861), .FEN(FEN[363]), .op(N861_t1) );
fim FAN_N867_0 ( .fault(fault), .net(N867), .FEN(FEN[364]), .op(N867_t0) );
fim FAN_N867_1 ( .fault(fault), .net(N867), .FEN(FEN[365]), .op(N867_t1) );
fim FAN_N870_0 ( .fault(fault), .net(N870), .FEN(FEN[366]), .op(N870_t0) );
fim FAN_N870_1 ( .fault(fault), .net(N870), .FEN(FEN[367]), .op(N870_t1) );
fim FAN_N870_2 ( .fault(fault), .net(N870), .FEN(FEN[368]), .op(N870_t2) );
fim FAN_N962_0 ( .fault(fault), .net(N962), .FEN(FEN[369]), .op(N962_t0) );
fim FAN_N962_1 ( .fault(fault), .net(N962), .FEN(FEN[370]), .op(N962_t1) );
fim FAN_N803_0 ( .fault(fault), .net(N803), .FEN(FEN[371]), .op(N803_t0) );
fim FAN_N803_1 ( .fault(fault), .net(N803), .FEN(FEN[372]), .op(N803_t1) );
fim FAN_N803_2 ( .fault(fault), .net(N803), .FEN(FEN[373]), .op(N803_t2) );
fim FAN_N803_3 ( .fault(fault), .net(N803), .FEN(FEN[374]), .op(N803_t3) );
fim FAN_N803_4 ( .fault(fault), .net(N803), .FEN(FEN[375]), .op(N803_t4) );
fim FAN_N803_5 ( .fault(fault), .net(N803), .FEN(FEN[376]), .op(N803_t5) );
fim FAN_N803_6 ( .fault(fault), .net(N803), .FEN(FEN[377]), .op(N803_t6) );
fim FAN_N803_7 ( .fault(fault), .net(N803), .FEN(FEN[378]), .op(N803_t7) );
fim FAN_N803_8 ( .fault(fault), .net(N803), .FEN(FEN[379]), .op(N803_t8) );
fim FAN_N803_9 ( .fault(fault), .net(N803), .FEN(FEN[380]), .op(N803_t9) );
fim FAN_N803_10 ( .fault(fault), .net(N803), .FEN(FEN[381]), .op(N803_t10) );
fim FAN_N803_11 ( .fault(fault), .net(N803), .FEN(FEN[382]), .op(N803_t11) );
fim FAN_N803_12 ( .fault(fault), .net(N803), .FEN(FEN[383]), .op(N803_t12) );
fim FAN_N803_13 ( .fault(fault), .net(N803), .FEN(FEN[384]), .op(N803_t13) );
fim FAN_N803_14 ( .fault(fault), .net(N803), .FEN(FEN[385]), .op(N803_t14) );
fim FAN_N803_15 ( .fault(fault), .net(N803), .FEN(FEN[386]), .op(N803_t15) );
fim FAN_N883_0 ( .fault(fault), .net(N883), .FEN(FEN[387]), .op(N883_t0) );
fim FAN_N883_1 ( .fault(fault), .net(N883), .FEN(FEN[388]), .op(N883_t1) );
fim FAN_N886_0 ( .fault(fault), .net(N886), .FEN(FEN[389]), .op(N886_t0) );
fim FAN_N886_1 ( .fault(fault), .net(N886), .FEN(FEN[390]), .op(N886_t1) );
fim FAN_N892_0 ( .fault(fault), .net(N892), .FEN(FEN[391]), .op(N892_t0) );
fim FAN_N892_1 ( .fault(fault), .net(N892), .FEN(FEN[392]), .op(N892_t1) );
fim FAN_N821_0 ( .fault(fault), .net(N821), .FEN(FEN[393]), .op(N821_t0) );
fim FAN_N821_1 ( .fault(fault), .net(N821), .FEN(FEN[394]), .op(N821_t1) );
fim FAN_N821_2 ( .fault(fault), .net(N821), .FEN(FEN[395]), .op(N821_t2) );
fim FAN_N896_0 ( .fault(fault), .net(N896), .FEN(FEN[396]), .op(N896_t0) );
fim FAN_N896_1 ( .fault(fault), .net(N896), .FEN(FEN[397]), .op(N896_t1) );
fim FAN_N896_2 ( .fault(fault), .net(N896), .FEN(FEN[398]), .op(N896_t2) );
fim FAN_N896_3 ( .fault(fault), .net(N896), .FEN(FEN[399]), .op(N896_t3) );
fim FAN_N896_4 ( .fault(fault), .net(N896), .FEN(FEN[400]), .op(N896_t4) );
fim FAN_N896_5 ( .fault(fault), .net(N896), .FEN(FEN[401]), .op(N896_t5) );
fim FAN_N896_6 ( .fault(fault), .net(N896), .FEN(FEN[402]), .op(N896_t6) );
fim FAN_N896_7 ( .fault(fault), .net(N896), .FEN(FEN[403]), .op(N896_t7) );
fim FAN_N896_8 ( .fault(fault), .net(N896), .FEN(FEN[404]), .op(N896_t8) );
fim FAN_N896_9 ( .fault(fault), .net(N896), .FEN(FEN[405]), .op(N896_t9) );
fim FAN_N896_10 ( .fault(fault), .net(N896), .FEN(FEN[406]), .op(N896_t10) );
fim FAN_N896_11 ( .fault(fault), .net(N896), .FEN(FEN[407]), .op(N896_t11) );
fim FAN_N896_12 ( .fault(fault), .net(N896), .FEN(FEN[408]), .op(N896_t12) );
fim FAN_N896_13 ( .fault(fault), .net(N896), .FEN(FEN[409]), .op(N896_t13) );
fim FAN_N896_14 ( .fault(fault), .net(N896), .FEN(FEN[410]), .op(N896_t14) );
fim FAN_N896_15 ( .fault(fault), .net(N896), .FEN(FEN[411]), .op(N896_t15) );
fim FAN_N829_0 ( .fault(fault), .net(N829), .FEN(FEN[412]), .op(N829_t0) );
fim FAN_N829_1 ( .fault(fault), .net(N829), .FEN(FEN[413]), .op(N829_t1) );
fim FAN_N917_0 ( .fault(fault), .net(N917), .FEN(FEN[414]), .op(N917_t0) );
fim FAN_N917_1 ( .fault(fault), .net(N917), .FEN(FEN[415]), .op(N917_t1) );
fim FAN_N965_0 ( .fault(fault), .net(N965), .FEN(FEN[416]), .op(N965_t0) );
fim FAN_N965_1 ( .fault(fault), .net(N965), .FEN(FEN[417]), .op(N965_t1) );
fim FAN_N920_0 ( .fault(fault), .net(N920), .FEN(FEN[418]), .op(N920_t0) );
fim FAN_N920_1 ( .fault(fault), .net(N920), .FEN(FEN[419]), .op(N920_t1) );
fim FAN_N923_0 ( .fault(fault), .net(N923), .FEN(FEN[420]), .op(N923_t0) );
fim FAN_N923_1 ( .fault(fault), .net(N923), .FEN(FEN[421]), .op(N923_t1) );
fim FAN_N938_0 ( .fault(fault), .net(N938), .FEN(FEN[422]), .op(N938_t0) );
fim FAN_N938_1 ( .fault(fault), .net(N938), .FEN(FEN[423]), .op(N938_t1) );
fim FAN_N941_0 ( .fault(fault), .net(N941), .FEN(FEN[424]), .op(N941_t0) );
fim FAN_N941_1 ( .fault(fault), .net(N941), .FEN(FEN[425]), .op(N941_t1) );
fim FAN_N944_0 ( .fault(fault), .net(N944), .FEN(FEN[426]), .op(N944_t0) );
fim FAN_N944_1 ( .fault(fault), .net(N944), .FEN(FEN[427]), .op(N944_t1) );
fim FAN_N947_0 ( .fault(fault), .net(N947), .FEN(FEN[428]), .op(N947_t0) );
fim FAN_N947_1 ( .fault(fault), .net(N947), .FEN(FEN[429]), .op(N947_t1) );
fim FAN_N950_0 ( .fault(fault), .net(N950), .FEN(FEN[430]), .op(N950_t0) );
fim FAN_N950_1 ( .fault(fault), .net(N950), .FEN(FEN[431]), .op(N950_t1) );
fim FAN_N702_0 ( .fault(fault), .net(N702), .FEN(FEN[432]), .op(N702_t0) );
fim FAN_N702_1 ( .fault(fault), .net(N702), .FEN(FEN[433]), .op(N702_t1) );
fim FAN_N702_2 ( .fault(fault), .net(N702), .FEN(FEN[434]), .op(N702_t2) );
fim FAN_N724_0 ( .fault(fault), .net(N724), .FEN(FEN[435]), .op(N724_t0) );
fim FAN_N724_1 ( .fault(fault), .net(N724), .FEN(FEN[436]), .op(N724_t1) );
fim FAN_N763_0 ( .fault(fault), .net(N763), .FEN(FEN[437]), .op(N763_t0) );
fim FAN_N763_1 ( .fault(fault), .net(N763), .FEN(FEN[438]), .op(N763_t1) );
fim FAN_N763_2 ( .fault(fault), .net(N763), .FEN(FEN[439]), .op(N763_t2) );
fim FAN_N763_3 ( .fault(fault), .net(N763), .FEN(FEN[440]), .op(N763_t3) );
fim FAN_N877_0 ( .fault(fault), .net(N877), .FEN(FEN[441]), .op(N877_t0) );
fim FAN_N877_1 ( .fault(fault), .net(N877), .FEN(FEN[442]), .op(N877_t1) );
fim FAN_N880_0 ( .fault(fault), .net(N880), .FEN(FEN[443]), .op(N880_t0) );
fim FAN_N880_1 ( .fault(fault), .net(N880), .FEN(FEN[444]), .op(N880_t1) );
fim FAN_N1117_0 ( .fault(fault), .net(N1117), .FEN(FEN[445]), .op(N1117_t0) );
fim FAN_N1117_1 ( .fault(fault), .net(N1117), .FEN(FEN[446]), .op(N1117_t1) );
fim FAN_N1117_2 ( .fault(fault), .net(N1117), .FEN(FEN[447]), .op(N1117_t2) );
fim FAN_N1117_3 ( .fault(fault), .net(N1117), .FEN(FEN[448]), .op(N1117_t3) );
fim FAN_N1117_4 ( .fault(fault), .net(N1117), .FEN(FEN[449]), .op(N1117_t4) );
fim FAN_N1117_5 ( .fault(fault), .net(N1117), .FEN(FEN[450]), .op(N1117_t5) );
fim FAN_N1117_6 ( .fault(fault), .net(N1117), .FEN(FEN[451]), .op(N1117_t6) );
fim FAN_N1117_7 ( .fault(fault), .net(N1117), .FEN(FEN[452]), .op(N1117_t7) );
fim FAN_N1117_8 ( .fault(fault), .net(N1117), .FEN(FEN[453]), .op(N1117_t8) );
fim FAN_N1117_9 ( .fault(fault), .net(N1117), .FEN(FEN[454]), .op(N1117_t9) );
fim FAN_N1117_10 ( .fault(fault), .net(N1117), .FEN(FEN[455]), .op(N1117_t10) );
fim FAN_N1117_11 ( .fault(fault), .net(N1117), .FEN(FEN[456]), .op(N1117_t11) );
fim FAN_N1117_12 ( .fault(fault), .net(N1117), .FEN(FEN[457]), .op(N1117_t12) );
fim FAN_N1117_13 ( .fault(fault), .net(N1117), .FEN(FEN[458]), .op(N1117_t13) );
fim FAN_N1117_14 ( .fault(fault), .net(N1117), .FEN(FEN[459]), .op(N1117_t14) );
fim FAN_N1117_15 ( .fault(fault), .net(N1117), .FEN(FEN[460]), .op(N1117_t15) );
fim FAN_N223_0 ( .fault(fault), .net(N223), .FEN(FEN[461]), .op(N223_t0) );
fim FAN_N223_1 ( .fault(fault), .net(N223), .FEN(FEN[462]), .op(N223_t1) );
fim FAN_N1202_0 ( .fault(fault), .net(N1202), .FEN(FEN[463]), .op(N1202_t0) );
fim FAN_N1202_1 ( .fault(fault), .net(N1202), .FEN(FEN[464]), .op(N1202_t1) );
fim FAN_N1202_2 ( .fault(fault), .net(N1202), .FEN(FEN[465]), .op(N1202_t2) );
fim FAN_N1202_3 ( .fault(fault), .net(N1202), .FEN(FEN[466]), .op(N1202_t3) );
fim FAN_N1202_4 ( .fault(fault), .net(N1202), .FEN(FEN[467]), .op(N1202_t4) );
fim FAN_N1202_5 ( .fault(fault), .net(N1202), .FEN(FEN[468]), .op(N1202_t5) );
fim FAN_N1202_6 ( .fault(fault), .net(N1202), .FEN(FEN[469]), .op(N1202_t6) );
fim FAN_N1202_7 ( .fault(fault), .net(N1202), .FEN(FEN[470]), .op(N1202_t7) );
fim FAN_N1202_8 ( .fault(fault), .net(N1202), .FEN(FEN[471]), .op(N1202_t8) );
fim FAN_N1202_9 ( .fault(fault), .net(N1202), .FEN(FEN[472]), .op(N1202_t9) );
fim FAN_N1202_10 ( .fault(fault), .net(N1202), .FEN(FEN[473]), .op(N1202_t10) );
fim FAN_N1202_11 ( .fault(fault), .net(N1202), .FEN(FEN[474]), .op(N1202_t11) );
fim FAN_N1202_12 ( .fault(fault), .net(N1202), .FEN(FEN[475]), .op(N1202_t12) );
fim FAN_N1202_13 ( .fault(fault), .net(N1202), .FEN(FEN[476]), .op(N1202_t13) );
fim FAN_N1202_14 ( .fault(fault), .net(N1202), .FEN(FEN[477]), .op(N1202_t14) );
fim FAN_N1202_15 ( .fault(fault), .net(N1202), .FEN(FEN[478]), .op(N1202_t15) );
fim FAN_N1264_0 ( .fault(fault), .net(N1264), .FEN(FEN[479]), .op(N1264_t0) );
fim FAN_N1264_1 ( .fault(fault), .net(N1264), .FEN(FEN[480]), .op(N1264_t1) );
fim FAN_N1340_0 ( .fault(fault), .net(N1340), .FEN(FEN[481]), .op(N1340_t0) );
fim FAN_N1340_1 ( .fault(fault), .net(N1340), .FEN(FEN[482]), .op(N1340_t1) );
fim FAN_N1268_0 ( .fault(fault), .net(N1268), .FEN(FEN[483]), .op(N1268_t0) );
fim FAN_N1268_1 ( .fault(fault), .net(N1268), .FEN(FEN[484]), .op(N1268_t1) );
fim FAN_N1493_0 ( .fault(fault), .net(N1493), .FEN(FEN[485]), .op(N1493_t0) );
fim FAN_N1493_1 ( .fault(fault), .net(N1493), .FEN(FEN[486]), .op(N1493_t1) );
fim FAN_N1499_0 ( .fault(fault), .net(N1499), .FEN(FEN[487]), .op(N1499_t0) );
fim FAN_N1499_1 ( .fault(fault), .net(N1499), .FEN(FEN[488]), .op(N1499_t1) );
fim FAN_N1273_0 ( .fault(fault), .net(N1273), .FEN(FEN[489]), .op(N1273_t0) );
fim FAN_N1273_1 ( .fault(fault), .net(N1273), .FEN(FEN[490]), .op(N1273_t1) );
fim FAN_N1276_0 ( .fault(fault), .net(N1276), .FEN(FEN[491]), .op(N1276_t0) );
fim FAN_N1276_1 ( .fault(fault), .net(N1276), .FEN(FEN[492]), .op(N1276_t1) );
fim FAN_N1325_0 ( .fault(fault), .net(N1325), .FEN(FEN[493]), .op(N1325_t0) );
fim FAN_N1325_1 ( .fault(fault), .net(N1325), .FEN(FEN[494]), .op(N1325_t1) );
fim FAN_N1279_0 ( .fault(fault), .net(N1279), .FEN(FEN[495]), .op(N1279_t0) );
fim FAN_N1279_1 ( .fault(fault), .net(N1279), .FEN(FEN[496]), .op(N1279_t1) );
fim FAN_N1302_0 ( .fault(fault), .net(N1302), .FEN(FEN[497]), .op(N1302_t0) );
fim FAN_N1302_1 ( .fault(fault), .net(N1302), .FEN(FEN[498]), .op(N1302_t1) );
fim FAN_N1302_2 ( .fault(fault), .net(N1302), .FEN(FEN[499]), .op(N1302_t2) );
fim FAN_N1496_0 ( .fault(fault), .net(N1496), .FEN(FEN[500]), .op(N1496_t0) );
fim FAN_N1496_1 ( .fault(fault), .net(N1496), .FEN(FEN[501]), .op(N1496_t1) );
fim FAN_N1502_0 ( .fault(fault), .net(N1502), .FEN(FEN[502]), .op(N1502_t0) );
fim FAN_N1502_1 ( .fault(fault), .net(N1502), .FEN(FEN[503]), .op(N1502_t1) );
fim FAN_N1328_0 ( .fault(fault), .net(N1328), .FEN(FEN[504]), .op(N1328_t0) );
fim FAN_N1328_1 ( .fault(fault), .net(N1328), .FEN(FEN[505]), .op(N1328_t1) );
fim FAN_N1334_0 ( .fault(fault), .net(N1334), .FEN(FEN[506]), .op(N1334_t0) );
fim FAN_N1334_1 ( .fault(fault), .net(N1334), .FEN(FEN[507]), .op(N1334_t1) );
fim FAN_N1331_0 ( .fault(fault), .net(N1331), .FEN(FEN[508]), .op(N1331_t0) );
fim FAN_N1331_1 ( .fault(fault), .net(N1331), .FEN(FEN[509]), .op(N1331_t1) );
fim FAN_N845_0 ( .fault(fault), .net(N845), .FEN(FEN[510]), .op(N845_t0) );
fim FAN_N845_1 ( .fault(fault), .net(N845), .FEN(FEN[511]), .op(N845_t1) );
fim FAN_N150_0 ( .fault(fault), .net(N150), .FEN(FEN[512]), .op(N150_t0) );
fim FAN_N150_1 ( .fault(fault), .net(N150), .FEN(FEN[513]), .op(N150_t1) );
fim FAN_N150_2 ( .fault(fault), .net(N150), .FEN(FEN[514]), .op(N150_t2) );
fim FAN_N150_3 ( .fault(fault), .net(N150), .FEN(FEN[515]), .op(N150_t3) );
fim FAN_N150_4 ( .fault(fault), .net(N150), .FEN(FEN[516]), .op(N150_t4) );
fim FAN_N150_5 ( .fault(fault), .net(N150), .FEN(FEN[517]), .op(N150_t5) );
fim FAN_N150_6 ( .fault(fault), .net(N150), .FEN(FEN[518]), .op(N150_t6) );
fim FAN_N150_7 ( .fault(fault), .net(N150), .FEN(FEN[519]), .op(N150_t7) );
fim FAN_N851_0 ( .fault(fault), .net(N851), .FEN(FEN[520]), .op(N851_t0) );
fim FAN_N851_1 ( .fault(fault), .net(N851), .FEN(FEN[521]), .op(N851_t1) );
fim FAN_N159_0 ( .fault(fault), .net(N159), .FEN(FEN[522]), .op(N159_t0) );
fim FAN_N159_1 ( .fault(fault), .net(N159), .FEN(FEN[523]), .op(N159_t1) );
fim FAN_N159_2 ( .fault(fault), .net(N159), .FEN(FEN[524]), .op(N159_t2) );
fim FAN_N159_3 ( .fault(fault), .net(N159), .FEN(FEN[525]), .op(N159_t3) );
fim FAN_N159_4 ( .fault(fault), .net(N159), .FEN(FEN[526]), .op(N159_t4) );
fim FAN_N159_5 ( .fault(fault), .net(N159), .FEN(FEN[527]), .op(N159_t5) );
fim FAN_N159_6 ( .fault(fault), .net(N159), .FEN(FEN[528]), .op(N159_t6) );
fim FAN_N159_7 ( .fault(fault), .net(N159), .FEN(FEN[529]), .op(N159_t7) );
fim FAN_N159_8 ( .fault(fault), .net(N159), .FEN(FEN[530]), .op(N159_t8) );
fim FAN_N858_0 ( .fault(fault), .net(N858), .FEN(FEN[531]), .op(N858_t0) );
fim FAN_N858_1 ( .fault(fault), .net(N858), .FEN(FEN[532]), .op(N858_t1) );
fim FAN_N864_0 ( .fault(fault), .net(N864), .FEN(FEN[533]), .op(N864_t0) );
fim FAN_N864_1 ( .fault(fault), .net(N864), .FEN(FEN[534]), .op(N864_t1) );
fim FAN_N283_0 ( .fault(fault), .net(N283), .FEN(FEN[535]), .op(N283_t0) );
fim FAN_N283_1 ( .fault(fault), .net(N283), .FEN(FEN[536]), .op(N283_t1) );
fim FAN_N283_2 ( .fault(fault), .net(N283), .FEN(FEN[537]), .op(N283_t2) );
fim FAN_N283_3 ( .fault(fault), .net(N283), .FEN(FEN[538]), .op(N283_t3) );
fim FAN_N283_4 ( .fault(fault), .net(N283), .FEN(FEN[539]), .op(N283_t4) );
fim FAN_N283_5 ( .fault(fault), .net(N283), .FEN(FEN[540]), .op(N283_t5) );
fim FAN_N283_6 ( .fault(fault), .net(N283), .FEN(FEN[541]), .op(N283_t6) );
fim FAN_N283_7 ( .fault(fault), .net(N283), .FEN(FEN[542]), .op(N283_t7) );
fim FAN_N283_8 ( .fault(fault), .net(N283), .FEN(FEN[543]), .op(N283_t8) );
fim FAN_N283_9 ( .fault(fault), .net(N283), .FEN(FEN[544]), .op(N283_t9) );
fim FAN_N1363_0 ( .fault(fault), .net(N1363), .FEN(FEN[545]), .op(N1363_t0) );
fim FAN_N1363_1 ( .fault(fault), .net(N1363), .FEN(FEN[546]), .op(N1363_t1) );
fim FAN_N1366_0 ( .fault(fault), .net(N1366), .FEN(FEN[547]), .op(N1366_t0) );
fim FAN_N1366_1 ( .fault(fault), .net(N1366), .FEN(FEN[548]), .op(N1366_t1) );
fim FAN_N1298_0 ( .fault(fault), .net(N1298), .FEN(FEN[549]), .op(N1298_t0) );
fim FAN_N1298_1 ( .fault(fault), .net(N1298), .FEN(FEN[550]), .op(N1298_t1) );
fim FAN_N1298_2 ( .fault(fault), .net(N1298), .FEN(FEN[551]), .op(N1298_t2) );
fim FAN_N1369_0 ( .fault(fault), .net(N1369), .FEN(FEN[552]), .op(N1369_t0) );
fim FAN_N1369_1 ( .fault(fault), .net(N1369), .FEN(FEN[553]), .op(N1369_t1) );
fim FAN_N1369_2 ( .fault(fault), .net(N1369), .FEN(FEN[554]), .op(N1369_t2) );
fim FAN_N1369_3 ( .fault(fault), .net(N1369), .FEN(FEN[555]), .op(N1369_t3) );
fim FAN_N1369_4 ( .fault(fault), .net(N1369), .FEN(FEN[556]), .op(N1369_t4) );
fim FAN_N1369_5 ( .fault(fault), .net(N1369), .FEN(FEN[557]), .op(N1369_t5) );
fim FAN_N1369_6 ( .fault(fault), .net(N1369), .FEN(FEN[558]), .op(N1369_t6) );
fim FAN_N1369_7 ( .fault(fault), .net(N1369), .FEN(FEN[559]), .op(N1369_t7) );
fim FAN_N1369_8 ( .fault(fault), .net(N1369), .FEN(FEN[560]), .op(N1369_t8) );
fim FAN_N1369_9 ( .fault(fault), .net(N1369), .FEN(FEN[561]), .op(N1369_t9) );
fim FAN_N1369_10 ( .fault(fault), .net(N1369), .FEN(FEN[562]), .op(N1369_t10) );
fim FAN_N1369_11 ( .fault(fault), .net(N1369), .FEN(FEN[563]), .op(N1369_t11) );
fim FAN_N1369_12 ( .fault(fault), .net(N1369), .FEN(FEN[564]), .op(N1369_t12) );
fim FAN_N1369_13 ( .fault(fault), .net(N1369), .FEN(FEN[565]), .op(N1369_t13) );
fim FAN_N1384_0 ( .fault(fault), .net(N1384), .FEN(FEN[566]), .op(N1384_t0) );
fim FAN_N1384_1 ( .fault(fault), .net(N1384), .FEN(FEN[567]), .op(N1384_t1) );
fim FAN_N1384_2 ( .fault(fault), .net(N1384), .FEN(FEN[568]), .op(N1384_t2) );
fim FAN_N1384_3 ( .fault(fault), .net(N1384), .FEN(FEN[569]), .op(N1384_t3) );
fim FAN_N1384_4 ( .fault(fault), .net(N1384), .FEN(FEN[570]), .op(N1384_t4) );
fim FAN_N1384_5 ( .fault(fault), .net(N1384), .FEN(FEN[571]), .op(N1384_t5) );
fim FAN_N1384_6 ( .fault(fault), .net(N1384), .FEN(FEN[572]), .op(N1384_t6) );
fim FAN_N1384_7 ( .fault(fault), .net(N1384), .FEN(FEN[573]), .op(N1384_t7) );
fim FAN_N1384_8 ( .fault(fault), .net(N1384), .FEN(FEN[574]), .op(N1384_t8) );
fim FAN_N1384_9 ( .fault(fault), .net(N1384), .FEN(FEN[575]), .op(N1384_t9) );
fim FAN_N1384_10 ( .fault(fault), .net(N1384), .FEN(FEN[576]), .op(N1384_t10) );
fim FAN_N1384_11 ( .fault(fault), .net(N1384), .FEN(FEN[577]), .op(N1384_t11) );
fim FAN_N1384_12 ( .fault(fault), .net(N1384), .FEN(FEN[578]), .op(N1384_t12) );
fim FAN_N1384_13 ( .fault(fault), .net(N1384), .FEN(FEN[579]), .op(N1384_t13) );
fim FAN_N1384_14 ( .fault(fault), .net(N1384), .FEN(FEN[580]), .op(N1384_t14) );
fim FAN_N1384_15 ( .fault(fault), .net(N1384), .FEN(FEN[581]), .op(N1384_t15) );
fim FAN_N1409_0 ( .fault(fault), .net(N1409), .FEN(FEN[582]), .op(N1409_t0) );
fim FAN_N1409_1 ( .fault(fault), .net(N1409), .FEN(FEN[583]), .op(N1409_t1) );
fim FAN_N1409_2 ( .fault(fault), .net(N1409), .FEN(FEN[584]), .op(N1409_t2) );
fim FAN_N1409_3 ( .fault(fault), .net(N1409), .FEN(FEN[585]), .op(N1409_t3) );
fim FAN_N1409_4 ( .fault(fault), .net(N1409), .FEN(FEN[586]), .op(N1409_t4) );
fim FAN_N1409_5 ( .fault(fault), .net(N1409), .FEN(FEN[587]), .op(N1409_t5) );
fim FAN_N1409_6 ( .fault(fault), .net(N1409), .FEN(FEN[588]), .op(N1409_t6) );
fim FAN_N1409_7 ( .fault(fault), .net(N1409), .FEN(FEN[589]), .op(N1409_t7) );
fim FAN_N1409_8 ( .fault(fault), .net(N1409), .FEN(FEN[590]), .op(N1409_t8) );
fim FAN_N1409_9 ( .fault(fault), .net(N1409), .FEN(FEN[591]), .op(N1409_t9) );
fim FAN_N1409_10 ( .fault(fault), .net(N1409), .FEN(FEN[592]), .op(N1409_t10) );
fim FAN_N1409_11 ( .fault(fault), .net(N1409), .FEN(FEN[593]), .op(N1409_t11) );
fim FAN_N1409_12 ( .fault(fault), .net(N1409), .FEN(FEN[594]), .op(N1409_t12) );
fim FAN_N1409_13 ( .fault(fault), .net(N1409), .FEN(FEN[595]), .op(N1409_t13) );
fim FAN_N1409_14 ( .fault(fault), .net(N1409), .FEN(FEN[596]), .op(N1409_t14) );
fim FAN_N1409_15 ( .fault(fault), .net(N1409), .FEN(FEN[597]), .op(N1409_t15) );
fim FAN_N1306_0 ( .fault(fault), .net(N1306), .FEN(FEN[598]), .op(N1306_t0) );
fim FAN_N1306_1 ( .fault(fault), .net(N1306), .FEN(FEN[599]), .op(N1306_t1) );
fim FAN_N1306_2 ( .fault(fault), .net(N1306), .FEN(FEN[600]), .op(N1306_t2) );
fim FAN_N1306_3 ( .fault(fault), .net(N1306), .FEN(FEN[601]), .op(N1306_t3) );
fim FAN_N1306_4 ( .fault(fault), .net(N1306), .FEN(FEN[602]), .op(N1306_t4) );
fim FAN_N1306_5 ( .fault(fault), .net(N1306), .FEN(FEN[603]), .op(N1306_t5) );
fim FAN_N1306_6 ( .fault(fault), .net(N1306), .FEN(FEN[604]), .op(N1306_t6) );
fim FAN_N1306_7 ( .fault(fault), .net(N1306), .FEN(FEN[605]), .op(N1306_t7) );
fim FAN_N1322_0 ( .fault(fault), .net(N1322), .FEN(FEN[606]), .op(N1322_t0) );
fim FAN_N1322_1 ( .fault(fault), .net(N1322), .FEN(FEN[607]), .op(N1322_t1) );
fim FAN_N1315_0 ( .fault(fault), .net(N1315), .FEN(FEN[608]), .op(N1315_t0) );
fim FAN_N1315_1 ( .fault(fault), .net(N1315), .FEN(FEN[609]), .op(N1315_t1) );
fim FAN_N1315_2 ( .fault(fault), .net(N1315), .FEN(FEN[610]), .op(N1315_t2) );
fim FAN_N1315_3 ( .fault(fault), .net(N1315), .FEN(FEN[611]), .op(N1315_t3) );
fim FAN_N1315_4 ( .fault(fault), .net(N1315), .FEN(FEN[612]), .op(N1315_t4) );
fim FAN_N1315_5 ( .fault(fault), .net(N1315), .FEN(FEN[613]), .op(N1315_t5) );
fim FAN_N1452_0 ( .fault(fault), .net(N1452), .FEN(FEN[614]), .op(N1452_t0) );
fim FAN_N1452_1 ( .fault(fault), .net(N1452), .FEN(FEN[615]), .op(N1452_t1) );
fim FAN_N1452_2 ( .fault(fault), .net(N1452), .FEN(FEN[616]), .op(N1452_t2) );
fim FAN_N1452_3 ( .fault(fault), .net(N1452), .FEN(FEN[617]), .op(N1452_t3) );
fim FAN_N1452_4 ( .fault(fault), .net(N1452), .FEN(FEN[618]), .op(N1452_t4) );
fim FAN_N1452_5 ( .fault(fault), .net(N1452), .FEN(FEN[619]), .op(N1452_t5) );
fim FAN_N1464_0 ( .fault(fault), .net(N1464), .FEN(FEN[620]), .op(N1464_t0) );
fim FAN_N1464_1 ( .fault(fault), .net(N1464), .FEN(FEN[621]), .op(N1464_t1) );
fim FAN_N1471_0 ( .fault(fault), .net(N1471), .FEN(FEN[622]), .op(N1471_t0) );
fim FAN_N1471_1 ( .fault(fault), .net(N1471), .FEN(FEN[623]), .op(N1471_t1) );
fim FAN_N1475_0 ( .fault(fault), .net(N1475), .FEN(FEN[624]), .op(N1475_t0) );
fim FAN_N1475_1 ( .fault(fault), .net(N1475), .FEN(FEN[625]), .op(N1475_t1) );
fim FAN_N1478_0 ( .fault(fault), .net(N1478), .FEN(FEN[626]), .op(N1478_t0) );
fim FAN_N1478_1 ( .fault(fault), .net(N1478), .FEN(FEN[627]), .op(N1478_t1) );
fim FAN_N1481_0 ( .fault(fault), .net(N1481), .FEN(FEN[628]), .op(N1481_t0) );
fim FAN_N1481_1 ( .fault(fault), .net(N1481), .FEN(FEN[629]), .op(N1481_t1) );
fim FAN_N1484_0 ( .fault(fault), .net(N1484), .FEN(FEN[630]), .op(N1484_t0) );
fim FAN_N1484_1 ( .fault(fault), .net(N1484), .FEN(FEN[631]), .op(N1484_t1) );
fim FAN_N1487_0 ( .fault(fault), .net(N1487), .FEN(FEN[632]), .op(N1487_t0) );
fim FAN_N1487_1 ( .fault(fault), .net(N1487), .FEN(FEN[633]), .op(N1487_t1) );
fim FAN_N1490_0 ( .fault(fault), .net(N1490), .FEN(FEN[634]), .op(N1490_t0) );
fim FAN_N1490_1 ( .fault(fault), .net(N1490), .FEN(FEN[635]), .op(N1490_t1) );
fim FAN_N1520_0 ( .fault(fault), .net(N1520), .FEN(FEN[636]), .op(N1520_t0) );
fim FAN_N1520_1 ( .fault(fault), .net(N1520), .FEN(FEN[637]), .op(N1520_t1) );
fim FAN_N1520_2 ( .fault(fault), .net(N1520), .FEN(FEN[638]), .op(N1520_t2) );
fim FAN_N294_0 ( .fault(fault), .net(N294), .FEN(FEN[639]), .op(N294_t0) );
fim FAN_N294_1 ( .fault(fault), .net(N294), .FEN(FEN[640]), .op(N294_t1) );
fim FAN_N294_2 ( .fault(fault), .net(N294), .FEN(FEN[641]), .op(N294_t2) );
fim FAN_N294_3 ( .fault(fault), .net(N294), .FEN(FEN[642]), .op(N294_t3) );
fim FAN_N294_4 ( .fault(fault), .net(N294), .FEN(FEN[643]), .op(N294_t4) );
fim FAN_N294_5 ( .fault(fault), .net(N294), .FEN(FEN[644]), .op(N294_t5) );
fim FAN_N294_6 ( .fault(fault), .net(N294), .FEN(FEN[645]), .op(N294_t6) );
fim FAN_N294_7 ( .fault(fault), .net(N294), .FEN(FEN[646]), .op(N294_t7) );
fim FAN_N303_0 ( .fault(fault), .net(N303), .FEN(FEN[647]), .op(N303_t0) );
fim FAN_N303_1 ( .fault(fault), .net(N303), .FEN(FEN[648]), .op(N303_t1) );
fim FAN_N303_2 ( .fault(fault), .net(N303), .FEN(FEN[649]), .op(N303_t2) );
fim FAN_N303_3 ( .fault(fault), .net(N303), .FEN(FEN[650]), .op(N303_t3) );
fim FAN_N303_4 ( .fault(fault), .net(N303), .FEN(FEN[651]), .op(N303_t4) );
fim FAN_N303_5 ( .fault(fault), .net(N303), .FEN(FEN[652]), .op(N303_t5) );
fim FAN_N303_6 ( .fault(fault), .net(N303), .FEN(FEN[653]), .op(N303_t6) );
fim FAN_N1667_0 ( .fault(fault), .net(N1667), .FEN(FEN[654]), .op(N1667_t0) );
fim FAN_N1667_1 ( .fault(fault), .net(N1667), .FEN(FEN[655]), .op(N1667_t1) );
fim FAN_N1670_0 ( .fault(fault), .net(N1670), .FEN(FEN[656]), .op(N1670_t0) );
fim FAN_N1670_1 ( .fault(fault), .net(N1670), .FEN(FEN[657]), .op(N1670_t1) );
fim FAN_N1197_0 ( .fault(fault), .net(N1197), .FEN(FEN[658]), .op(N1197_t0) );
fim FAN_N1197_1 ( .fault(fault), .net(N1197), .FEN(FEN[659]), .op(N1197_t1) );
fim FAN_N1197_2 ( .fault(fault), .net(N1197), .FEN(FEN[660]), .op(N1197_t2) );
fim FAN_N1197_3 ( .fault(fault), .net(N1197), .FEN(FEN[661]), .op(N1197_t3) );
fim FAN_N1219_0 ( .fault(fault), .net(N1219), .FEN(FEN[662]), .op(N1219_t0) );
fim FAN_N1219_1 ( .fault(fault), .net(N1219), .FEN(FEN[663]), .op(N1219_t1) );
fim FAN_N1219_2 ( .fault(fault), .net(N1219), .FEN(FEN[664]), .op(N1219_t2) );
fim FAN_N1219_3 ( .fault(fault), .net(N1219), .FEN(FEN[665]), .op(N1219_t3) );
fim FAN_N1562_0 ( .fault(fault), .net(N1562), .FEN(FEN[666]), .op(N1562_t0) );
fim FAN_N1562_1 ( .fault(fault), .net(N1562), .FEN(FEN[667]), .op(N1562_t1) );
fim FAN_N1562_2 ( .fault(fault), .net(N1562), .FEN(FEN[668]), .op(N1562_t2) );
fim FAN_N1562_3 ( .fault(fault), .net(N1562), .FEN(FEN[669]), .op(N1562_t3) );
fim FAN_N1562_4 ( .fault(fault), .net(N1562), .FEN(FEN[670]), .op(N1562_t4) );
fim FAN_N1562_5 ( .fault(fault), .net(N1562), .FEN(FEN[671]), .op(N1562_t5) );
fim FAN_N1562_6 ( .fault(fault), .net(N1562), .FEN(FEN[672]), .op(N1562_t6) );
fim FAN_N1562_7 ( .fault(fault), .net(N1562), .FEN(FEN[673]), .op(N1562_t7) );
fim FAN_N1562_8 ( .fault(fault), .net(N1562), .FEN(FEN[674]), .op(N1562_t8) );
fim FAN_N1562_9 ( .fault(fault), .net(N1562), .FEN(FEN[675]), .op(N1562_t9) );
fim FAN_N1562_10 ( .fault(fault), .net(N1562), .FEN(FEN[676]), .op(N1562_t10) );
fim FAN_N1562_11 ( .fault(fault), .net(N1562), .FEN(FEN[677]), .op(N1562_t11) );
fim FAN_N1562_12 ( .fault(fault), .net(N1562), .FEN(FEN[678]), .op(N1562_t12) );
fim FAN_N1562_13 ( .fault(fault), .net(N1562), .FEN(FEN[679]), .op(N1562_t13) );
fim FAN_N1562_14 ( .fault(fault), .net(N1562), .FEN(FEN[680]), .op(N1562_t14) );
fim FAN_N1562_15 ( .fault(fault), .net(N1562), .FEN(FEN[681]), .op(N1562_t15) );
fim FAN_N1933_0 ( .fault(fault), .net(N1933), .FEN(FEN[682]), .op(N1933_t0) );
fim FAN_N1933_1 ( .fault(fault), .net(N1933), .FEN(FEN[683]), .op(N1933_t1) );
fim FAN_N1936_0 ( .fault(fault), .net(N1936), .FEN(FEN[684]), .op(N1936_t0) );
fim FAN_N1936_1 ( .fault(fault), .net(N1936), .FEN(FEN[685]), .op(N1936_t1) );
fim FAN_N1738_0 ( .fault(fault), .net(N1738), .FEN(FEN[686]), .op(N1738_t0) );
fim FAN_N1738_1 ( .fault(fault), .net(N1738), .FEN(FEN[687]), .op(N1738_t1) );
fim FAN_N1738_2 ( .fault(fault), .net(N1738), .FEN(FEN[688]), .op(N1738_t2) );
fim FAN_N1738_3 ( .fault(fault), .net(N1738), .FEN(FEN[689]), .op(N1738_t3) );
fim FAN_N1738_4 ( .fault(fault), .net(N1738), .FEN(FEN[690]), .op(N1738_t4) );
fim FAN_N1738_5 ( .fault(fault), .net(N1738), .FEN(FEN[691]), .op(N1738_t5) );
fim FAN_N1738_6 ( .fault(fault), .net(N1738), .FEN(FEN[692]), .op(N1738_t6) );
fim FAN_N1738_7 ( .fault(fault), .net(N1738), .FEN(FEN[693]), .op(N1738_t7) );
fim FAN_N1747_0 ( .fault(fault), .net(N1747), .FEN(FEN[694]), .op(N1747_t0) );
fim FAN_N1747_1 ( .fault(fault), .net(N1747), .FEN(FEN[695]), .op(N1747_t1) );
fim FAN_N1747_2 ( .fault(fault), .net(N1747), .FEN(FEN[696]), .op(N1747_t2) );
fim FAN_N1747_3 ( .fault(fault), .net(N1747), .FEN(FEN[697]), .op(N1747_t3) );
fim FAN_N1747_4 ( .fault(fault), .net(N1747), .FEN(FEN[698]), .op(N1747_t4) );
fim FAN_N1747_5 ( .fault(fault), .net(N1747), .FEN(FEN[699]), .op(N1747_t5) );
fim FAN_N1747_6 ( .fault(fault), .net(N1747), .FEN(FEN[700]), .op(N1747_t6) );
fim FAN_N1747_7 ( .fault(fault), .net(N1747), .FEN(FEN[701]), .op(N1747_t7) );
fim FAN_N1722_0 ( .fault(fault), .net(N1722), .FEN(FEN[702]), .op(N1722_t0) );
fim FAN_N1722_1 ( .fault(fault), .net(N1722), .FEN(FEN[703]), .op(N1722_t1) );
fim FAN_N1761_0 ( .fault(fault), .net(N1761), .FEN(FEN[704]), .op(N1761_t0) );
fim FAN_N1761_1 ( .fault(fault), .net(N1761), .FEN(FEN[705]), .op(N1761_t1) );
fim FAN_N1756_0 ( .fault(fault), .net(N1756), .FEN(FEN[706]), .op(N1756_t0) );
fim FAN_N1756_1 ( .fault(fault), .net(N1756), .FEN(FEN[707]), .op(N1756_t1) );
fim FAN_N1756_2 ( .fault(fault), .net(N1756), .FEN(FEN[708]), .op(N1756_t2) );
fim FAN_N1756_3 ( .fault(fault), .net(N1756), .FEN(FEN[709]), .op(N1756_t3) );
fim FAN_N1358_0 ( .fault(fault), .net(N1358), .FEN(FEN[710]), .op(N1358_t0) );
fim FAN_N1358_1 ( .fault(fault), .net(N1358), .FEN(FEN[711]), .op(N1358_t1) );
fim FAN_N1358_2 ( .fault(fault), .net(N1358), .FEN(FEN[712]), .op(N1358_t2) );
fim FAN_N1358_3 ( .fault(fault), .net(N1358), .FEN(FEN[713]), .op(N1358_t3) );
fim FAN_N1812_0 ( .fault(fault), .net(N1812), .FEN(FEN[714]), .op(N1812_t0) );
fim FAN_N1812_1 ( .fault(fault), .net(N1812), .FEN(FEN[715]), .op(N1812_t1) );
fim FAN_N1809_0 ( .fault(fault), .net(N1809), .FEN(FEN[716]), .op(N1809_t0) );
fim FAN_N1809_1 ( .fault(fault), .net(N1809), .FEN(FEN[717]), .op(N1809_t1) );
fim FAN_N1353_0 ( .fault(fault), .net(N1353), .FEN(FEN[718]), .op(N1353_t0) );
fim FAN_N1353_1 ( .fault(fault), .net(N1353), .FEN(FEN[719]), .op(N1353_t1) );
fim FAN_N1353_2 ( .fault(fault), .net(N1353), .FEN(FEN[720]), .op(N1353_t2) );
fim FAN_N1353_3 ( .fault(fault), .net(N1353), .FEN(FEN[721]), .op(N1353_t3) );
fim FAN_N1806_0 ( .fault(fault), .net(N1806), .FEN(FEN[722]), .op(N1806_t0) );
fim FAN_N1806_1 ( .fault(fault), .net(N1806), .FEN(FEN[723]), .op(N1806_t1) );
fim FAN_N1803_0 ( .fault(fault), .net(N1803), .FEN(FEN[724]), .op(N1803_t0) );
fim FAN_N1803_1 ( .fault(fault), .net(N1803), .FEN(FEN[725]), .op(N1803_t1) );
fim FAN_N1815_0 ( .fault(fault), .net(N1815), .FEN(FEN[726]), .op(N1815_t0) );
fim FAN_N1815_1 ( .fault(fault), .net(N1815), .FEN(FEN[727]), .op(N1815_t1) );
fim FAN_N1818_0 ( .fault(fault), .net(N1818), .FEN(FEN[728]), .op(N1818_t0) );
fim FAN_N1818_1 ( .fault(fault), .net(N1818), .FEN(FEN[729]), .op(N1818_t1) );
fim FAN_N1821_0 ( .fault(fault), .net(N1821), .FEN(FEN[730]), .op(N1821_t0) );
fim FAN_N1821_1 ( .fault(fault), .net(N1821), .FEN(FEN[731]), .op(N1821_t1) );
fim FAN_N1833_0 ( .fault(fault), .net(N1833), .FEN(FEN[732]), .op(N1833_t0) );
fim FAN_N1833_1 ( .fault(fault), .net(N1833), .FEN(FEN[733]), .op(N1833_t1) );
fim FAN_N1833_2 ( .fault(fault), .net(N1833), .FEN(FEN[734]), .op(N1833_t2) );
fim FAN_N1833_3 ( .fault(fault), .net(N1833), .FEN(FEN[735]), .op(N1833_t3) );
fim FAN_N1833_4 ( .fault(fault), .net(N1833), .FEN(FEN[736]), .op(N1833_t4) );
fim FAN_N1833_5 ( .fault(fault), .net(N1833), .FEN(FEN[737]), .op(N1833_t5) );
fim FAN_N1833_6 ( .fault(fault), .net(N1833), .FEN(FEN[738]), .op(N1833_t6) );
fim FAN_N1833_7 ( .fault(fault), .net(N1833), .FEN(FEN[739]), .op(N1833_t7) );
fim FAN_N1824_0 ( .fault(fault), .net(N1824), .FEN(FEN[740]), .op(N1824_t0) );
fim FAN_N1824_1 ( .fault(fault), .net(N1824), .FEN(FEN[741]), .op(N1824_t1) );
fim FAN_N1824_2 ( .fault(fault), .net(N1824), .FEN(FEN[742]), .op(N1824_t2) );
fim FAN_N1824_3 ( .fault(fault), .net(N1824), .FEN(FEN[743]), .op(N1824_t3) );
fim FAN_N1824_4 ( .fault(fault), .net(N1824), .FEN(FEN[744]), .op(N1824_t4) );
fim FAN_N1824_5 ( .fault(fault), .net(N1824), .FEN(FEN[745]), .op(N1824_t5) );
fim FAN_N1824_6 ( .fault(fault), .net(N1824), .FEN(FEN[746]), .op(N1824_t6) );
fim FAN_N1824_7 ( .fault(fault), .net(N1824), .FEN(FEN[747]), .op(N1824_t7) );
fim FAN_N1917_0 ( .fault(fault), .net(N1917), .FEN(FEN[748]), .op(N1917_t0) );
fim FAN_N1917_1 ( .fault(fault), .net(N1917), .FEN(FEN[749]), .op(N1917_t1) );
fim FAN_N1917_2 ( .fault(fault), .net(N1917), .FEN(FEN[750]), .op(N1917_t2) );
fim FAN_N1917_3 ( .fault(fault), .net(N1917), .FEN(FEN[751]), .op(N1917_t3) );
fim FAN_N1930_0 ( .fault(fault), .net(N1930), .FEN(FEN[752]), .op(N1930_t0) );
fim FAN_N1930_1 ( .fault(fault), .net(N1930), .FEN(FEN[753]), .op(N1930_t1) );
fim FAN_N350_0 ( .fault(fault), .net(N350), .FEN(FEN[754]), .op(N350_t0) );
fim FAN_N350_1 ( .fault(fault), .net(N350), .FEN(FEN[755]), .op(N350_t1) );
fim FAN_N1715_0 ( .fault(fault), .net(N1715), .FEN(FEN[756]), .op(N1715_t0) );
fim FAN_N1715_1 ( .fault(fault), .net(N1715), .FEN(FEN[757]), .op(N1715_t1) );
fim FAN_N1718_0 ( .fault(fault), .net(N1718), .FEN(FEN[758]), .op(N1718_t0) );
fim FAN_N1718_1 ( .fault(fault), .net(N1718), .FEN(FEN[759]), .op(N1718_t1) );
fim FAN_N2057_0 ( .fault(fault), .net(N2057), .FEN(FEN[760]), .op(N2057_t0) );
fim FAN_N2057_1 ( .fault(fault), .net(N2057), .FEN(FEN[761]), .op(N2057_t1) );
fim FAN_N2057_2 ( .fault(fault), .net(N2057), .FEN(FEN[762]), .op(N2057_t2) );
fim FAN_N2057_3 ( .fault(fault), .net(N2057), .FEN(FEN[763]), .op(N2057_t3) );
fim FAN_N2057_4 ( .fault(fault), .net(N2057), .FEN(FEN[764]), .op(N2057_t4) );
fim FAN_N2057_5 ( .fault(fault), .net(N2057), .FEN(FEN[765]), .op(N2057_t5) );
fim FAN_N2057_6 ( .fault(fault), .net(N2057), .FEN(FEN[766]), .op(N2057_t6) );
fim FAN_N2057_7 ( .fault(fault), .net(N2057), .FEN(FEN[767]), .op(N2057_t7) );
fim FAN_N274_0 ( .fault(fault), .net(N274), .FEN(FEN[768]), .op(N274_t0) );
fim FAN_N274_1 ( .fault(fault), .net(N274), .FEN(FEN[769]), .op(N274_t1) );
fim FAN_N274_2 ( .fault(fault), .net(N274), .FEN(FEN[770]), .op(N274_t2) );
fim FAN_N274_3 ( .fault(fault), .net(N274), .FEN(FEN[771]), .op(N274_t3) );
fim FAN_N274_4 ( .fault(fault), .net(N274), .FEN(FEN[772]), .op(N274_t4) );
fim FAN_N274_5 ( .fault(fault), .net(N274), .FEN(FEN[773]), .op(N274_t5) );
fim FAN_N274_6 ( .fault(fault), .net(N274), .FEN(FEN[774]), .op(N274_t6) );
fim FAN_N274_7 ( .fault(fault), .net(N274), .FEN(FEN[775]), .op(N274_t7) );
fim FAN_N2052_0 ( .fault(fault), .net(N2052), .FEN(FEN[776]), .op(N2052_t0) );
fim FAN_N2052_1 ( .fault(fault), .net(N2052), .FEN(FEN[777]), .op(N2052_t1) );
fim FAN_N2052_2 ( .fault(fault), .net(N2052), .FEN(FEN[778]), .op(N2052_t2) );
fim FAN_N2052_3 ( .fault(fault), .net(N2052), .FEN(FEN[779]), .op(N2052_t3) );
fim FAN_N2043_0 ( .fault(fault), .net(N2043), .FEN(FEN[780]), .op(N2043_t0) );
fim FAN_N2043_1 ( .fault(fault), .net(N2043), .FEN(FEN[781]), .op(N2043_t1) );
fim FAN_N2043_2 ( .fault(fault), .net(N2043), .FEN(FEN[782]), .op(N2043_t2) );
fim FAN_N2043_3 ( .fault(fault), .net(N2043), .FEN(FEN[783]), .op(N2043_t3) );
fim FAN_N2043_4 ( .fault(fault), .net(N2043), .FEN(FEN[784]), .op(N2043_t4) );
fim FAN_N2043_5 ( .fault(fault), .net(N2043), .FEN(FEN[785]), .op(N2043_t5) );
fim FAN_N2043_6 ( .fault(fault), .net(N2043), .FEN(FEN[786]), .op(N2043_t6) );
fim FAN_N2043_7 ( .fault(fault), .net(N2043), .FEN(FEN[787]), .op(N2043_t7) );
fim FAN_N2038_0 ( .fault(fault), .net(N2038), .FEN(FEN[788]), .op(N2038_t0) );
fim FAN_N2038_1 ( .fault(fault), .net(N2038), .FEN(FEN[789]), .op(N2038_t1) );
fim FAN_N2038_2 ( .fault(fault), .net(N2038), .FEN(FEN[790]), .op(N2038_t2) );
fim FAN_N2038_3 ( .fault(fault), .net(N2038), .FEN(FEN[791]), .op(N2038_t3) );
fim FAN_N2313_0 ( .fault(fault), .net(N2313), .FEN(FEN[792]), .op(N2313_t0) );
fim FAN_N2313_1 ( .fault(fault), .net(N2313), .FEN(FEN[793]), .op(N2313_t1) );
fim FAN_N2316_0 ( .fault(fault), .net(N2316), .FEN(FEN[794]), .op(N2316_t0) );
fim FAN_N2316_1 ( .fault(fault), .net(N2316), .FEN(FEN[795]), .op(N2316_t1) );
fim FAN_N2319_0 ( .fault(fault), .net(N2319), .FEN(FEN[796]), .op(N2319_t0) );
fim FAN_N2319_1 ( .fault(fault), .net(N2319), .FEN(FEN[797]), .op(N2319_t1) );
fim FAN_N2322_0 ( .fault(fault), .net(N2322), .FEN(FEN[798]), .op(N2322_t0) );
fim FAN_N2322_1 ( .fault(fault), .net(N2322), .FEN(FEN[799]), .op(N2322_t1) );
fim FAN_N2325_0 ( .fault(fault), .net(N2325), .FEN(FEN[800]), .op(N2325_t0) );
fim FAN_N2325_1 ( .fault(fault), .net(N2325), .FEN(FEN[801]), .op(N2325_t1) );
fim FAN_N2328_0 ( .fault(fault), .net(N2328), .FEN(FEN[802]), .op(N2328_t0) );
fim FAN_N2328_1 ( .fault(fault), .net(N2328), .FEN(FEN[803]), .op(N2328_t1) );
fim FAN_N2331_0 ( .fault(fault), .net(N2331), .FEN(FEN[804]), .op(N2331_t0) );
fim FAN_N2331_1 ( .fault(fault), .net(N2331), .FEN(FEN[805]), .op(N2331_t1) );
fim FAN_N2334_0 ( .fault(fault), .net(N2334), .FEN(FEN[806]), .op(N2334_t0) );
fim FAN_N2334_1 ( .fault(fault), .net(N2334), .FEN(FEN[807]), .op(N2334_t1) );
fim FAN_N2175_0 ( .fault(fault), .net(N2175), .FEN(FEN[808]), .op(N2175_t0) );
fim FAN_N2175_1 ( .fault(fault), .net(N2175), .FEN(FEN[809]), .op(N2175_t1) );
fim FAN_N2185_0 ( .fault(fault), .net(N2185), .FEN(FEN[810]), .op(N2185_t0) );
fim FAN_N2185_1 ( .fault(fault), .net(N2185), .FEN(FEN[811]), .op(N2185_t1) );
fim FAN_N2188_0 ( .fault(fault), .net(N2188), .FEN(FEN[812]), .op(N2188_t0) );
fim FAN_N2188_1 ( .fault(fault), .net(N2188), .FEN(FEN[813]), .op(N2188_t1) );
fim FAN_N2191_0 ( .fault(fault), .net(N2191), .FEN(FEN[814]), .op(N2191_t0) );
fim FAN_N2191_1 ( .fault(fault), .net(N2191), .FEN(FEN[815]), .op(N2191_t1) );
fim FAN_N2194_0 ( .fault(fault), .net(N2194), .FEN(FEN[816]), .op(N2194_t0) );
fim FAN_N2194_1 ( .fault(fault), .net(N2194), .FEN(FEN[817]), .op(N2194_t1) );
fim FAN_N2197_0 ( .fault(fault), .net(N2197), .FEN(FEN[818]), .op(N2197_t0) );
fim FAN_N2197_1 ( .fault(fault), .net(N2197), .FEN(FEN[819]), .op(N2197_t1) );
fim FAN_N2200_0 ( .fault(fault), .net(N2200), .FEN(FEN[820]), .op(N2200_t0) );
fim FAN_N2200_1 ( .fault(fault), .net(N2200), .FEN(FEN[821]), .op(N2200_t1) );
fim FAN_N2203_0 ( .fault(fault), .net(N2203), .FEN(FEN[822]), .op(N2203_t0) );
fim FAN_N2203_1 ( .fault(fault), .net(N2203), .FEN(FEN[823]), .op(N2203_t1) );
fim FAN_N2206_0 ( .fault(fault), .net(N2206), .FEN(FEN[824]), .op(N2206_t0) );
fim FAN_N2206_1 ( .fault(fault), .net(N2206), .FEN(FEN[825]), .op(N2206_t1) );
fim FAN_N2212_0 ( .fault(fault), .net(N2212), .FEN(FEN[826]), .op(N2212_t0) );
fim FAN_N2212_1 ( .fault(fault), .net(N2212), .FEN(FEN[827]), .op(N2212_t1) );
fim FAN_N2212_2 ( .fault(fault), .net(N2212), .FEN(FEN[828]), .op(N2212_t2) );
fim FAN_N2212_3 ( .fault(fault), .net(N2212), .FEN(FEN[829]), .op(N2212_t3) );
fim FAN_N2212_4 ( .fault(fault), .net(N2212), .FEN(FEN[830]), .op(N2212_t4) );
fim FAN_N2212_5 ( .fault(fault), .net(N2212), .FEN(FEN[831]), .op(N2212_t5) );
fim FAN_N2212_6 ( .fault(fault), .net(N2212), .FEN(FEN[832]), .op(N2212_t6) );
fim FAN_N2212_7 ( .fault(fault), .net(N2212), .FEN(FEN[833]), .op(N2212_t7) );
fim FAN_N2221_0 ( .fault(fault), .net(N2221), .FEN(FEN[834]), .op(N2221_t0) );
fim FAN_N2221_1 ( .fault(fault), .net(N2221), .FEN(FEN[835]), .op(N2221_t1) );
fim FAN_N2221_2 ( .fault(fault), .net(N2221), .FEN(FEN[836]), .op(N2221_t2) );
fim FAN_N2221_3 ( .fault(fault), .net(N2221), .FEN(FEN[837]), .op(N2221_t3) );
fim FAN_N2221_4 ( .fault(fault), .net(N2221), .FEN(FEN[838]), .op(N2221_t4) );
fim FAN_N2221_5 ( .fault(fault), .net(N2221), .FEN(FEN[839]), .op(N2221_t5) );
fim FAN_N2221_6 ( .fault(fault), .net(N2221), .FEN(FEN[840]), .op(N2221_t6) );
fim FAN_N2221_7 ( .fault(fault), .net(N2221), .FEN(FEN[841]), .op(N2221_t7) );
fim FAN_N2270_0 ( .fault(fault), .net(N2270), .FEN(FEN[842]), .op(N2270_t0) );
fim FAN_N2270_1 ( .fault(fault), .net(N2270), .FEN(FEN[843]), .op(N2270_t1) );
fim FAN_N1870_0 ( .fault(fault), .net(N1870), .FEN(FEN[844]), .op(N1870_t0) );
fim FAN_N1870_1 ( .fault(fault), .net(N1870), .FEN(FEN[845]), .op(N1870_t1) );
fim FAN_N2068_0 ( .fault(fault), .net(N2068), .FEN(FEN[846]), .op(N2068_t0) );
fim FAN_N2068_1 ( .fault(fault), .net(N2068), .FEN(FEN[847]), .op(N2068_t1) );
fim FAN_N2277_0 ( .fault(fault), .net(N2277), .FEN(FEN[848]), .op(N2277_t0) );
fim FAN_N2277_1 ( .fault(fault), .net(N2277), .FEN(FEN[849]), .op(N2277_t1) );
fim FAN_N1880_0 ( .fault(fault), .net(N1880), .FEN(FEN[850]), .op(N1880_t0) );
fim FAN_N1880_1 ( .fault(fault), .net(N1880), .FEN(FEN[851]), .op(N1880_t1) );
fim FAN_N2078_0 ( .fault(fault), .net(N2078), .FEN(FEN[852]), .op(N2078_t0) );
fim FAN_N2078_1 ( .fault(fault), .net(N2078), .FEN(FEN[853]), .op(N2078_t1) );
fim FAN_N2282_0 ( .fault(fault), .net(N2282), .FEN(FEN[854]), .op(N2282_t0) );
fim FAN_N2282_1 ( .fault(fault), .net(N2282), .FEN(FEN[855]), .op(N2282_t1) );
fim FAN_N1885_0 ( .fault(fault), .net(N1885), .FEN(FEN[856]), .op(N1885_t0) );
fim FAN_N1885_1 ( .fault(fault), .net(N1885), .FEN(FEN[857]), .op(N1885_t1) );
fim FAN_N2083_0 ( .fault(fault), .net(N2083), .FEN(FEN[858]), .op(N2083_t0) );
fim FAN_N2083_1 ( .fault(fault), .net(N2083), .FEN(FEN[859]), .op(N2083_t1) );
fim FAN_N2287_0 ( .fault(fault), .net(N2287), .FEN(FEN[860]), .op(N2287_t0) );
fim FAN_N2287_1 ( .fault(fault), .net(N2287), .FEN(FEN[861]), .op(N2287_t1) );
fim FAN_N1890_0 ( .fault(fault), .net(N1890), .FEN(FEN[862]), .op(N1890_t0) );
fim FAN_N1890_1 ( .fault(fault), .net(N1890), .FEN(FEN[863]), .op(N1890_t1) );
fim FAN_N2088_0 ( .fault(fault), .net(N2088), .FEN(FEN[864]), .op(N2088_t0) );
fim FAN_N2088_1 ( .fault(fault), .net(N2088), .FEN(FEN[865]), .op(N2088_t1) );
fim FAN_N2294_0 ( .fault(fault), .net(N2294), .FEN(FEN[866]), .op(N2294_t0) );
fim FAN_N2294_1 ( .fault(fault), .net(N2294), .FEN(FEN[867]), .op(N2294_t1) );
fim FAN_N1900_0 ( .fault(fault), .net(N1900), .FEN(FEN[868]), .op(N1900_t0) );
fim FAN_N1900_1 ( .fault(fault), .net(N1900), .FEN(FEN[869]), .op(N1900_t1) );
fim FAN_N2098_0 ( .fault(fault), .net(N2098), .FEN(FEN[870]), .op(N2098_t0) );
fim FAN_N2098_1 ( .fault(fault), .net(N2098), .FEN(FEN[871]), .op(N2098_t1) );
fim FAN_N2299_0 ( .fault(fault), .net(N2299), .FEN(FEN[872]), .op(N2299_t0) );
fim FAN_N2299_1 ( .fault(fault), .net(N2299), .FEN(FEN[873]), .op(N2299_t1) );
fim FAN_N1905_0 ( .fault(fault), .net(N1905), .FEN(FEN[874]), .op(N1905_t0) );
fim FAN_N1905_1 ( .fault(fault), .net(N1905), .FEN(FEN[875]), .op(N1905_t1) );
fim FAN_N2103_0 ( .fault(fault), .net(N2103), .FEN(FEN[876]), .op(N2103_t0) );
fim FAN_N2103_1 ( .fault(fault), .net(N2103), .FEN(FEN[877]), .op(N2103_t1) );
fim FAN_N2304_0 ( .fault(fault), .net(N2304), .FEN(FEN[878]), .op(N2304_t0) );
fim FAN_N2304_1 ( .fault(fault), .net(N2304), .FEN(FEN[879]), .op(N2304_t1) );
fim FAN_N2158_0 ( .fault(fault), .net(N2158), .FEN(FEN[880]), .op(N2158_t0) );
fim FAN_N2158_1 ( .fault(fault), .net(N2158), .FEN(FEN[881]), .op(N2158_t1) );
fim FAN_N2158_2 ( .fault(fault), .net(N2158), .FEN(FEN[882]), .op(N2158_t2) );
fim FAN_N2158_3 ( .fault(fault), .net(N2158), .FEN(FEN[883]), .op(N2158_t3) );
fim FAN_N2158_4 ( .fault(fault), .net(N2158), .FEN(FEN[884]), .op(N2158_t4) );
fim FAN_N2158_5 ( .fault(fault), .net(N2158), .FEN(FEN[885]), .op(N2158_t5) );
fim FAN_N2158_6 ( .fault(fault), .net(N2158), .FEN(FEN[886]), .op(N2158_t6) );
fim FAN_N2158_7 ( .fault(fault), .net(N2158), .FEN(FEN[887]), .op(N2158_t7) );
fim FAN_N2158_8 ( .fault(fault), .net(N2158), .FEN(FEN[888]), .op(N2158_t8) );
fim FAN_N2158_9 ( .fault(fault), .net(N2158), .FEN(FEN[889]), .op(N2158_t9) );
fim FAN_N2158_10 ( .fault(fault), .net(N2158), .FEN(FEN[890]), .op(N2158_t10) );
fim FAN_N2158_11 ( .fault(fault), .net(N2158), .FEN(FEN[891]), .op(N2158_t11) );
fim FAN_N2158_12 ( .fault(fault), .net(N2158), .FEN(FEN[892]), .op(N2158_t12) );
fim FAN_N2158_13 ( .fault(fault), .net(N2158), .FEN(FEN[893]), .op(N2158_t13) );
fim FAN_N2158_14 ( .fault(fault), .net(N2158), .FEN(FEN[894]), .op(N2158_t14) );
fim FAN_N2158_15 ( .fault(fault), .net(N2158), .FEN(FEN[895]), .op(N2158_t15) );
fim FAN_N2376_0 ( .fault(fault), .net(N2376), .FEN(FEN[896]), .op(N2376_t0) );
fim FAN_N2376_1 ( .fault(fault), .net(N2376), .FEN(FEN[897]), .op(N2376_t1) );
fim FAN_N1983_0 ( .fault(fault), .net(N1983), .FEN(FEN[898]), .op(N1983_t0) );
fim FAN_N1983_1 ( .fault(fault), .net(N1983), .FEN(FEN[899]), .op(N1983_t1) );
fim FAN_N2379_0 ( .fault(fault), .net(N2379), .FEN(FEN[900]), .op(N2379_t0) );
fim FAN_N2379_1 ( .fault(fault), .net(N2379), .FEN(FEN[901]), .op(N2379_t1) );
fim FAN_N2471_0 ( .fault(fault), .net(N2471), .FEN(FEN[902]), .op(N2471_t0) );
fim FAN_N2471_1 ( .fault(fault), .net(N2471), .FEN(FEN[903]), .op(N2471_t1) );
fim FAN_N2488_0 ( .fault(fault), .net(N2488), .FEN(FEN[904]), .op(N2488_t0) );
fim FAN_N2488_1 ( .fault(fault), .net(N2488), .FEN(FEN[905]), .op(N2488_t1) );
fim FAN_N2488_2 ( .fault(fault), .net(N2488), .FEN(FEN[906]), .op(N2488_t2) );
fim FAN_N2488_3 ( .fault(fault), .net(N2488), .FEN(FEN[907]), .op(N2488_t3) );
fim FAN_N2488_4 ( .fault(fault), .net(N2488), .FEN(FEN[908]), .op(N2488_t4) );
fim FAN_N2488_5 ( .fault(fault), .net(N2488), .FEN(FEN[909]), .op(N2488_t5) );
fim FAN_N2488_6 ( .fault(fault), .net(N2488), .FEN(FEN[910]), .op(N2488_t6) );
fim FAN_N2488_7 ( .fault(fault), .net(N2488), .FEN(FEN[911]), .op(N2488_t7) );
fim FAN_N2497_0 ( .fault(fault), .net(N2497), .FEN(FEN[912]), .op(N2497_t0) );
fim FAN_N2497_1 ( .fault(fault), .net(N2497), .FEN(FEN[913]), .op(N2497_t1) );
fim FAN_N2497_2 ( .fault(fault), .net(N2497), .FEN(FEN[914]), .op(N2497_t2) );
fim FAN_N2497_3 ( .fault(fault), .net(N2497), .FEN(FEN[915]), .op(N2497_t3) );
fim FAN_N2497_4 ( .fault(fault), .net(N2497), .FEN(FEN[916]), .op(N2497_t4) );
fim FAN_N2497_5 ( .fault(fault), .net(N2497), .FEN(FEN[917]), .op(N2497_t5) );
fim FAN_N2497_6 ( .fault(fault), .net(N2497), .FEN(FEN[918]), .op(N2497_t6) );
fim FAN_N2497_7 ( .fault(fault), .net(N2497), .FEN(FEN[919]), .op(N2497_t7) );
fim FAN_N2506_0 ( .fault(fault), .net(N2506), .FEN(FEN[920]), .op(N2506_t0) );
fim FAN_N2506_1 ( .fault(fault), .net(N2506), .FEN(FEN[921]), .op(N2506_t1) );
fim FAN_N2506_2 ( .fault(fault), .net(N2506), .FEN(FEN[922]), .op(N2506_t2) );
fim FAN_N2506_3 ( .fault(fault), .net(N2506), .FEN(FEN[923]), .op(N2506_t3) );
fim FAN_N2506_4 ( .fault(fault), .net(N2506), .FEN(FEN[924]), .op(N2506_t4) );
fim FAN_N2506_5 ( .fault(fault), .net(N2506), .FEN(FEN[925]), .op(N2506_t5) );
fim FAN_N2506_6 ( .fault(fault), .net(N2506), .FEN(FEN[926]), .op(N2506_t6) );
fim FAN_N2506_7 ( .fault(fault), .net(N2506), .FEN(FEN[927]), .op(N2506_t7) );
fim FAN_N2515_0 ( .fault(fault), .net(N2515), .FEN(FEN[928]), .op(N2515_t0) );
fim FAN_N2515_1 ( .fault(fault), .net(N2515), .FEN(FEN[929]), .op(N2515_t1) );
fim FAN_N2515_2 ( .fault(fault), .net(N2515), .FEN(FEN[930]), .op(N2515_t2) );
fim FAN_N2515_3 ( .fault(fault), .net(N2515), .FEN(FEN[931]), .op(N2515_t3) );
fim FAN_N2515_4 ( .fault(fault), .net(N2515), .FEN(FEN[932]), .op(N2515_t4) );
fim FAN_N2515_5 ( .fault(fault), .net(N2515), .FEN(FEN[933]), .op(N2515_t5) );
fim FAN_N2515_6 ( .fault(fault), .net(N2515), .FEN(FEN[934]), .op(N2515_t6) );
fim FAN_N2515_7 ( .fault(fault), .net(N2515), .FEN(FEN[935]), .op(N2515_t7) );
fim FAN_N2524_0 ( .fault(fault), .net(N2524), .FEN(FEN[936]), .op(N2524_t0) );
fim FAN_N2524_1 ( .fault(fault), .net(N2524), .FEN(FEN[937]), .op(N2524_t1) );
fim FAN_N2524_2 ( .fault(fault), .net(N2524), .FEN(FEN[938]), .op(N2524_t2) );
fim FAN_N2524_3 ( .fault(fault), .net(N2524), .FEN(FEN[939]), .op(N2524_t3) );
fim FAN_N2524_4 ( .fault(fault), .net(N2524), .FEN(FEN[940]), .op(N2524_t4) );
fim FAN_N2524_5 ( .fault(fault), .net(N2524), .FEN(FEN[941]), .op(N2524_t5) );
fim FAN_N2524_6 ( .fault(fault), .net(N2524), .FEN(FEN[942]), .op(N2524_t6) );
fim FAN_N2524_7 ( .fault(fault), .net(N2524), .FEN(FEN[943]), .op(N2524_t7) );
fim FAN_N2533_0 ( .fault(fault), .net(N2533), .FEN(FEN[944]), .op(N2533_t0) );
fim FAN_N2533_1 ( .fault(fault), .net(N2533), .FEN(FEN[945]), .op(N2533_t1) );
fim FAN_N2533_2 ( .fault(fault), .net(N2533), .FEN(FEN[946]), .op(N2533_t2) );
fim FAN_N2533_3 ( .fault(fault), .net(N2533), .FEN(FEN[947]), .op(N2533_t3) );
fim FAN_N2533_4 ( .fault(fault), .net(N2533), .FEN(FEN[948]), .op(N2533_t4) );
fim FAN_N2533_5 ( .fault(fault), .net(N2533), .FEN(FEN[949]), .op(N2533_t5) );
fim FAN_N2533_6 ( .fault(fault), .net(N2533), .FEN(FEN[950]), .op(N2533_t6) );
fim FAN_N2533_7 ( .fault(fault), .net(N2533), .FEN(FEN[951]), .op(N2533_t7) );
fim FAN_N2542_0 ( .fault(fault), .net(N2542), .FEN(FEN[952]), .op(N2542_t0) );
fim FAN_N2542_1 ( .fault(fault), .net(N2542), .FEN(FEN[953]), .op(N2542_t1) );
fim FAN_N2542_2 ( .fault(fault), .net(N2542), .FEN(FEN[954]), .op(N2542_t2) );
fim FAN_N2542_3 ( .fault(fault), .net(N2542), .FEN(FEN[955]), .op(N2542_t3) );
fim FAN_N2542_4 ( .fault(fault), .net(N2542), .FEN(FEN[956]), .op(N2542_t4) );
fim FAN_N2542_5 ( .fault(fault), .net(N2542), .FEN(FEN[957]), .op(N2542_t5) );
fim FAN_N2542_6 ( .fault(fault), .net(N2542), .FEN(FEN[958]), .op(N2542_t6) );
fim FAN_N2542_7 ( .fault(fault), .net(N2542), .FEN(FEN[959]), .op(N2542_t7) );
fim FAN_N2551_0 ( .fault(fault), .net(N2551), .FEN(FEN[960]), .op(N2551_t0) );
fim FAN_N2551_1 ( .fault(fault), .net(N2551), .FEN(FEN[961]), .op(N2551_t1) );
fim FAN_N2551_2 ( .fault(fault), .net(N2551), .FEN(FEN[962]), .op(N2551_t2) );
fim FAN_N2551_3 ( .fault(fault), .net(N2551), .FEN(FEN[963]), .op(N2551_t3) );
fim FAN_N2551_4 ( .fault(fault), .net(N2551), .FEN(FEN[964]), .op(N2551_t4) );
fim FAN_N2551_5 ( .fault(fault), .net(N2551), .FEN(FEN[965]), .op(N2551_t5) );
fim FAN_N2551_6 ( .fault(fault), .net(N2551), .FEN(FEN[966]), .op(N2551_t6) );
fim FAN_N2551_7 ( .fault(fault), .net(N2551), .FEN(FEN[967]), .op(N2551_t7) );
fim FAN_N2560_0 ( .fault(fault), .net(N2560), .FEN(FEN[968]), .op(N2560_t0) );
fim FAN_N2560_1 ( .fault(fault), .net(N2560), .FEN(FEN[969]), .op(N2560_t1) );
fim FAN_N2560_2 ( .fault(fault), .net(N2560), .FEN(FEN[970]), .op(N2560_t2) );
fim FAN_N2560_3 ( .fault(fault), .net(N2560), .FEN(FEN[971]), .op(N2560_t3) );
fim FAN_N2560_4 ( .fault(fault), .net(N2560), .FEN(FEN[972]), .op(N2560_t4) );
fim FAN_N2560_5 ( .fault(fault), .net(N2560), .FEN(FEN[973]), .op(N2560_t5) );
fim FAN_N2560_6 ( .fault(fault), .net(N2560), .FEN(FEN[974]), .op(N2560_t6) );
fim FAN_N2560_7 ( .fault(fault), .net(N2560), .FEN(FEN[975]), .op(N2560_t7) );
fim FAN_N2569_0 ( .fault(fault), .net(N2569), .FEN(FEN[976]), .op(N2569_t0) );
fim FAN_N2569_1 ( .fault(fault), .net(N2569), .FEN(FEN[977]), .op(N2569_t1) );
fim FAN_N2569_2 ( .fault(fault), .net(N2569), .FEN(FEN[978]), .op(N2569_t2) );
fim FAN_N2569_3 ( .fault(fault), .net(N2569), .FEN(FEN[979]), .op(N2569_t3) );
fim FAN_N2569_4 ( .fault(fault), .net(N2569), .FEN(FEN[980]), .op(N2569_t4) );
fim FAN_N2569_5 ( .fault(fault), .net(N2569), .FEN(FEN[981]), .op(N2569_t5) );
fim FAN_N2569_6 ( .fault(fault), .net(N2569), .FEN(FEN[982]), .op(N2569_t6) );
fim FAN_N2569_7 ( .fault(fault), .net(N2569), .FEN(FEN[983]), .op(N2569_t7) );
fim FAN_N2578_0 ( .fault(fault), .net(N2578), .FEN(FEN[984]), .op(N2578_t0) );
fim FAN_N2578_1 ( .fault(fault), .net(N2578), .FEN(FEN[985]), .op(N2578_t1) );
fim FAN_N2578_2 ( .fault(fault), .net(N2578), .FEN(FEN[986]), .op(N2578_t2) );
fim FAN_N2578_3 ( .fault(fault), .net(N2578), .FEN(FEN[987]), .op(N2578_t3) );
fim FAN_N2578_4 ( .fault(fault), .net(N2578), .FEN(FEN[988]), .op(N2578_t4) );
fim FAN_N2578_5 ( .fault(fault), .net(N2578), .FEN(FEN[989]), .op(N2578_t5) );
fim FAN_N2578_6 ( .fault(fault), .net(N2578), .FEN(FEN[990]), .op(N2578_t6) );
fim FAN_N2578_7 ( .fault(fault), .net(N2578), .FEN(FEN[991]), .op(N2578_t7) );
fim FAN_N2587_0 ( .fault(fault), .net(N2587), .FEN(FEN[992]), .op(N2587_t0) );
fim FAN_N2587_1 ( .fault(fault), .net(N2587), .FEN(FEN[993]), .op(N2587_t1) );
fim FAN_N2587_2 ( .fault(fault), .net(N2587), .FEN(FEN[994]), .op(N2587_t2) );
fim FAN_N2587_3 ( .fault(fault), .net(N2587), .FEN(FEN[995]), .op(N2587_t3) );
fim FAN_N2587_4 ( .fault(fault), .net(N2587), .FEN(FEN[996]), .op(N2587_t4) );
fim FAN_N2587_5 ( .fault(fault), .net(N2587), .FEN(FEN[997]), .op(N2587_t5) );
fim FAN_N2587_6 ( .fault(fault), .net(N2587), .FEN(FEN[998]), .op(N2587_t6) );
fim FAN_N2587_7 ( .fault(fault), .net(N2587), .FEN(FEN[999]), .op(N2587_t7) );
fim FAN_N2596_0 ( .fault(fault), .net(N2596), .FEN(FEN[1000]), .op(N2596_t0) );
fim FAN_N2596_1 ( .fault(fault), .net(N2596), .FEN(FEN[1001]), .op(N2596_t1) );
fim FAN_N2596_2 ( .fault(fault), .net(N2596), .FEN(FEN[1002]), .op(N2596_t2) );
fim FAN_N2596_3 ( .fault(fault), .net(N2596), .FEN(FEN[1003]), .op(N2596_t3) );
fim FAN_N2596_4 ( .fault(fault), .net(N2596), .FEN(FEN[1004]), .op(N2596_t4) );
fim FAN_N2596_5 ( .fault(fault), .net(N2596), .FEN(FEN[1005]), .op(N2596_t5) );
fim FAN_N2596_6 ( .fault(fault), .net(N2596), .FEN(FEN[1006]), .op(N2596_t6) );
fim FAN_N2596_7 ( .fault(fault), .net(N2596), .FEN(FEN[1007]), .op(N2596_t7) );
fim FAN_N2605_0 ( .fault(fault), .net(N2605), .FEN(FEN[1008]), .op(N2605_t0) );
fim FAN_N2605_1 ( .fault(fault), .net(N2605), .FEN(FEN[1009]), .op(N2605_t1) );
fim FAN_N2605_2 ( .fault(fault), .net(N2605), .FEN(FEN[1010]), .op(N2605_t2) );
fim FAN_N2605_3 ( .fault(fault), .net(N2605), .FEN(FEN[1011]), .op(N2605_t3) );
fim FAN_N2605_4 ( .fault(fault), .net(N2605), .FEN(FEN[1012]), .op(N2605_t4) );
fim FAN_N2605_5 ( .fault(fault), .net(N2605), .FEN(FEN[1013]), .op(N2605_t5) );
fim FAN_N2605_6 ( .fault(fault), .net(N2605), .FEN(FEN[1014]), .op(N2605_t6) );
fim FAN_N2605_7 ( .fault(fault), .net(N2605), .FEN(FEN[1015]), .op(N2605_t7) );
fim FAN_N2614_0 ( .fault(fault), .net(N2614), .FEN(FEN[1016]), .op(N2614_t0) );
fim FAN_N2614_1 ( .fault(fault), .net(N2614), .FEN(FEN[1017]), .op(N2614_t1) );
fim FAN_N2614_2 ( .fault(fault), .net(N2614), .FEN(FEN[1018]), .op(N2614_t2) );
fim FAN_N2614_3 ( .fault(fault), .net(N2614), .FEN(FEN[1019]), .op(N2614_t3) );
fim FAN_N2614_4 ( .fault(fault), .net(N2614), .FEN(FEN[1020]), .op(N2614_t4) );
fim FAN_N2614_5 ( .fault(fault), .net(N2614), .FEN(FEN[1021]), .op(N2614_t5) );
fim FAN_N2614_6 ( .fault(fault), .net(N2614), .FEN(FEN[1022]), .op(N2614_t6) );
fim FAN_N2614_7 ( .fault(fault), .net(N2614), .FEN(FEN[1023]), .op(N2614_t7) );
fim FAN_N2623_0 ( .fault(fault), .net(N2623), .FEN(FEN[1024]), .op(N2623_t0) );
fim FAN_N2623_1 ( .fault(fault), .net(N2623), .FEN(FEN[1025]), .op(N2623_t1) );
fim FAN_N2623_2 ( .fault(fault), .net(N2623), .FEN(FEN[1026]), .op(N2623_t2) );
fim FAN_N2623_3 ( .fault(fault), .net(N2623), .FEN(FEN[1027]), .op(N2623_t3) );
fim FAN_N2623_4 ( .fault(fault), .net(N2623), .FEN(FEN[1028]), .op(N2623_t4) );
fim FAN_N2623_5 ( .fault(fault), .net(N2623), .FEN(FEN[1029]), .op(N2623_t5) );
fim FAN_N2623_6 ( .fault(fault), .net(N2623), .FEN(FEN[1030]), .op(N2623_t6) );
fim FAN_N2623_7 ( .fault(fault), .net(N2623), .FEN(FEN[1031]), .op(N2623_t7) );
fim FAN_N2656_0 ( .fault(fault), .net(N2656), .FEN(FEN[1032]), .op(N2656_t0) );
fim FAN_N2656_1 ( .fault(fault), .net(N2656), .FEN(FEN[1033]), .op(N2656_t1) );
fim FAN_N2652_0 ( .fault(fault), .net(N2652), .FEN(FEN[1034]), .op(N2652_t0) );
fim FAN_N2652_1 ( .fault(fault), .net(N2652), .FEN(FEN[1035]), .op(N2652_t1) );
fim FAN_N2652_2 ( .fault(fault), .net(N2652), .FEN(FEN[1036]), .op(N2652_t2) );
fim FAN_N2659_0 ( .fault(fault), .net(N2659), .FEN(FEN[1037]), .op(N2659_t0) );
fim FAN_N2659_1 ( .fault(fault), .net(N2659), .FEN(FEN[1038]), .op(N2659_t1) );
fim FAN_N2670_0 ( .fault(fault), .net(N2670), .FEN(FEN[1039]), .op(N2670_t0) );
fim FAN_N2670_1 ( .fault(fault), .net(N2670), .FEN(FEN[1040]), .op(N2670_t1) );
fim FAN_N2666_0 ( .fault(fault), .net(N2666), .FEN(FEN[1041]), .op(N2666_t0) );
fim FAN_N2666_1 ( .fault(fault), .net(N2666), .FEN(FEN[1042]), .op(N2666_t1) );
fim FAN_N2666_2 ( .fault(fault), .net(N2666), .FEN(FEN[1043]), .op(N2666_t2) );
fim FAN_N2681_0 ( .fault(fault), .net(N2681), .FEN(FEN[1044]), .op(N2681_t0) );
fim FAN_N2681_1 ( .fault(fault), .net(N2681), .FEN(FEN[1045]), .op(N2681_t1) );
fim FAN_N2677_0 ( .fault(fault), .net(N2677), .FEN(FEN[1046]), .op(N2677_t0) );
fim FAN_N2677_1 ( .fault(fault), .net(N2677), .FEN(FEN[1047]), .op(N2677_t1) );
fim FAN_N2677_2 ( .fault(fault), .net(N2677), .FEN(FEN[1048]), .op(N2677_t2) );
fim FAN_N2692_0 ( .fault(fault), .net(N2692), .FEN(FEN[1049]), .op(N2692_t0) );
fim FAN_N2692_1 ( .fault(fault), .net(N2692), .FEN(FEN[1050]), .op(N2692_t1) );
fim FAN_N2692_2 ( .fault(fault), .net(N2692), .FEN(FEN[1051]), .op(N2692_t2) );
fim FAN_N2692_3 ( .fault(fault), .net(N2692), .FEN(FEN[1052]), .op(N2692_t3) );
fim FAN_N2688_0 ( .fault(fault), .net(N2688), .FEN(FEN[1053]), .op(N2688_t0) );
fim FAN_N2688_1 ( .fault(fault), .net(N2688), .FEN(FEN[1054]), .op(N2688_t1) );
fim FAN_N2688_2 ( .fault(fault), .net(N2688), .FEN(FEN[1055]), .op(N2688_t2) );
fim FAN_N2697_0 ( .fault(fault), .net(N2697), .FEN(FEN[1056]), .op(N2697_t0) );
fim FAN_N2697_1 ( .fault(fault), .net(N2697), .FEN(FEN[1057]), .op(N2697_t1) );
fim FAN_N2697_2 ( .fault(fault), .net(N2697), .FEN(FEN[1058]), .op(N2697_t2) );
fim FAN_N2697_3 ( .fault(fault), .net(N2697), .FEN(FEN[1059]), .op(N2697_t3) );
fim FAN_N2710_0 ( .fault(fault), .net(N2710), .FEN(FEN[1060]), .op(N2710_t0) );
fim FAN_N2710_1 ( .fault(fault), .net(N2710), .FEN(FEN[1061]), .op(N2710_t1) );
fim FAN_N2710_2 ( .fault(fault), .net(N2710), .FEN(FEN[1062]), .op(N2710_t2) );
fim FAN_N2710_3 ( .fault(fault), .net(N2710), .FEN(FEN[1063]), .op(N2710_t3) );
fim FAN_N2706_0 ( .fault(fault), .net(N2706), .FEN(FEN[1064]), .op(N2706_t0) );
fim FAN_N2706_1 ( .fault(fault), .net(N2706), .FEN(FEN[1065]), .op(N2706_t1) );
fim FAN_N2706_2 ( .fault(fault), .net(N2706), .FEN(FEN[1066]), .op(N2706_t2) );
fim FAN_N2723_0 ( .fault(fault), .net(N2723), .FEN(FEN[1067]), .op(N2723_t0) );
fim FAN_N2723_1 ( .fault(fault), .net(N2723), .FEN(FEN[1068]), .op(N2723_t1) );
fim FAN_N2723_2 ( .fault(fault), .net(N2723), .FEN(FEN[1069]), .op(N2723_t2) );
fim FAN_N2723_3 ( .fault(fault), .net(N2723), .FEN(FEN[1070]), .op(N2723_t3) );
fim FAN_N2719_0 ( .fault(fault), .net(N2719), .FEN(FEN[1071]), .op(N2719_t0) );
fim FAN_N2719_1 ( .fault(fault), .net(N2719), .FEN(FEN[1072]), .op(N2719_t1) );
fim FAN_N2719_2 ( .fault(fault), .net(N2719), .FEN(FEN[1073]), .op(N2719_t2) );
fim FAN_N1909_0 ( .fault(fault), .net(N1909), .FEN(FEN[1074]), .op(N1909_t0) );
fim FAN_N1909_1 ( .fault(fault), .net(N1909), .FEN(FEN[1075]), .op(N1909_t1) );
fim FAN_N2648_0 ( .fault(fault), .net(N2648), .FEN(FEN[1076]), .op(N2648_t0) );
fim FAN_N2648_1 ( .fault(fault), .net(N2648), .FEN(FEN[1077]), .op(N2648_t1) );
fim FAN_N2648_2 ( .fault(fault), .net(N2648), .FEN(FEN[1078]), .op(N2648_t2) );
fim FAN_N1913_0 ( .fault(fault), .net(N1913), .FEN(FEN[1079]), .op(N1913_t0) );
fim FAN_N1913_1 ( .fault(fault), .net(N1913), .FEN(FEN[1080]), .op(N1913_t1) );
fim FAN_N1913_2 ( .fault(fault), .net(N1913), .FEN(FEN[1081]), .op(N1913_t2) );
fim FAN_N2662_0 ( .fault(fault), .net(N2662), .FEN(FEN[1082]), .op(N2662_t0) );
fim FAN_N2662_1 ( .fault(fault), .net(N2662), .FEN(FEN[1083]), .op(N2662_t1) );
fim FAN_N2662_2 ( .fault(fault), .net(N2662), .FEN(FEN[1084]), .op(N2662_t2) );
fim FAN_N2673_0 ( .fault(fault), .net(N2673), .FEN(FEN[1085]), .op(N2673_t0) );
fim FAN_N2673_1 ( .fault(fault), .net(N2673), .FEN(FEN[1086]), .op(N2673_t1) );
fim FAN_N2673_2 ( .fault(fault), .net(N2673), .FEN(FEN[1087]), .op(N2673_t2) );
fim FAN_N2684_0 ( .fault(fault), .net(N2684), .FEN(FEN[1088]), .op(N2684_t0) );
fim FAN_N2684_1 ( .fault(fault), .net(N2684), .FEN(FEN[1089]), .op(N2684_t1) );
fim FAN_N2684_2 ( .fault(fault), .net(N2684), .FEN(FEN[1090]), .op(N2684_t2) );
fim FAN_N1922_0 ( .fault(fault), .net(N1922), .FEN(FEN[1091]), .op(N1922_t0) );
fim FAN_N1922_1 ( .fault(fault), .net(N1922), .FEN(FEN[1092]), .op(N1922_t1) );
fim FAN_N1922_2 ( .fault(fault), .net(N1922), .FEN(FEN[1093]), .op(N1922_t2) );
fim FAN_N2702_0 ( .fault(fault), .net(N2702), .FEN(FEN[1094]), .op(N2702_t0) );
fim FAN_N2702_1 ( .fault(fault), .net(N2702), .FEN(FEN[1095]), .op(N2702_t1) );
fim FAN_N2702_2 ( .fault(fault), .net(N2702), .FEN(FEN[1096]), .op(N2702_t2) );
fim FAN_N2715_0 ( .fault(fault), .net(N2715), .FEN(FEN[1097]), .op(N2715_t0) );
fim FAN_N2715_1 ( .fault(fault), .net(N2715), .FEN(FEN[1098]), .op(N2715_t1) );
fim FAN_N2715_2 ( .fault(fault), .net(N2715), .FEN(FEN[1099]), .op(N2715_t2) );
fim FAN_N143_0 ( .fault(fault), .net(N143), .FEN(FEN[1100]), .op(N143_t0) );
fim FAN_N143_1 ( .fault(fault), .net(N143), .FEN(FEN[1101]), .op(N143_t1) );
fim FAN_N143_2 ( .fault(fault), .net(N143), .FEN(FEN[1102]), .op(N143_t2) );
fim FAN_N143_3 ( .fault(fault), .net(N143), .FEN(FEN[1103]), .op(N143_t3) );
fim FAN_N143_4 ( .fault(fault), .net(N143), .FEN(FEN[1104]), .op(N143_t4) );
fim FAN_N143_5 ( .fault(fault), .net(N143), .FEN(FEN[1105]), .op(N143_t5) );
fim FAN_N137_0 ( .fault(fault), .net(N137), .FEN(FEN[1106]), .op(N137_t0) );
fim FAN_N137_1 ( .fault(fault), .net(N137), .FEN(FEN[1107]), .op(N137_t1) );
fim FAN_N137_2 ( .fault(fault), .net(N137), .FEN(FEN[1108]), .op(N137_t2) );
fim FAN_N137_3 ( .fault(fault), .net(N137), .FEN(FEN[1109]), .op(N137_t3) );
fim FAN_N137_4 ( .fault(fault), .net(N137), .FEN(FEN[1110]), .op(N137_t4) );
fim FAN_N132_0 ( .fault(fault), .net(N132), .FEN(FEN[1111]), .op(N132_t0) );
fim FAN_N132_1 ( .fault(fault), .net(N132), .FEN(FEN[1112]), .op(N132_t1) );
fim FAN_N132_2 ( .fault(fault), .net(N132), .FEN(FEN[1113]), .op(N132_t2) );
fim FAN_N132_3 ( .fault(fault), .net(N132), .FEN(FEN[1114]), .op(N132_t3) );
fim FAN_N128_0 ( .fault(fault), .net(N128), .FEN(FEN[1115]), .op(N128_t0) );
fim FAN_N128_1 ( .fault(fault), .net(N128), .FEN(FEN[1116]), .op(N128_t1) );
fim FAN_N128_2 ( .fault(fault), .net(N128), .FEN(FEN[1117]), .op(N128_t2) );
fim FAN_N125_0 ( .fault(fault), .net(N125), .FEN(FEN[1118]), .op(N125_t0) );
fim FAN_N125_1 ( .fault(fault), .net(N125), .FEN(FEN[1119]), .op(N125_t1) );
fim FAN_N311_0 ( .fault(fault), .net(N311), .FEN(FEN[1120]), .op(N311_t0) );
fim FAN_N311_1 ( .fault(fault), .net(N311), .FEN(FEN[1121]), .op(N311_t1) );
fim FAN_N311_2 ( .fault(fault), .net(N311), .FEN(FEN[1122]), .op(N311_t2) );
fim FAN_N311_3 ( .fault(fault), .net(N311), .FEN(FEN[1123]), .op(N311_t3) );
fim FAN_N311_4 ( .fault(fault), .net(N311), .FEN(FEN[1124]), .op(N311_t4) );
fim FAN_N317_0 ( .fault(fault), .net(N317), .FEN(FEN[1125]), .op(N317_t0) );
fim FAN_N317_1 ( .fault(fault), .net(N317), .FEN(FEN[1126]), .op(N317_t1) );
fim FAN_N317_2 ( .fault(fault), .net(N317), .FEN(FEN[1127]), .op(N317_t2) );
fim FAN_N317_3 ( .fault(fault), .net(N317), .FEN(FEN[1128]), .op(N317_t3) );
fim FAN_N322_0 ( .fault(fault), .net(N322), .FEN(FEN[1129]), .op(N322_t0) );
fim FAN_N322_1 ( .fault(fault), .net(N322), .FEN(FEN[1130]), .op(N322_t1) );
fim FAN_N322_2 ( .fault(fault), .net(N322), .FEN(FEN[1131]), .op(N322_t2) );
fim FAN_N326_0 ( .fault(fault), .net(N326), .FEN(FEN[1132]), .op(N326_t0) );
fim FAN_N326_1 ( .fault(fault), .net(N326), .FEN(FEN[1133]), .op(N326_t1) );
fim FAN_N2977_0 ( .fault(fault), .net(N2977), .FEN(FEN[1134]), .op(N2977_t0) );
fim FAN_N2977_1 ( .fault(fault), .net(N2977), .FEN(FEN[1135]), .op(N2977_t1) );
fim FAN_N2973_0 ( .fault(fault), .net(N2973), .FEN(FEN[1136]), .op(N2973_t0) );
fim FAN_N2973_1 ( .fault(fault), .net(N2973), .FEN(FEN[1137]), .op(N2973_t1) );
fim FAN_N2973_2 ( .fault(fault), .net(N2973), .FEN(FEN[1138]), .op(N2973_t2) );
fim FAN_N3112_0 ( .fault(fault), .net(N3112), .FEN(FEN[1139]), .op(N3112_t0) );
fim FAN_N3112_1 ( .fault(fault), .net(N3112), .FEN(FEN[1140]), .op(N3112_t1) );
fim FAN_N3115_0 ( .fault(fault), .net(N3115), .FEN(FEN[1141]), .op(N3115_t0) );
fim FAN_N3115_1 ( .fault(fault), .net(N3115), .FEN(FEN[1142]), .op(N3115_t1) );
fim FAN_N3119_0 ( .fault(fault), .net(N3119), .FEN(FEN[1143]), .op(N3119_t0) );
fim FAN_N3119_1 ( .fault(fault), .net(N3119), .FEN(FEN[1144]), .op(N3119_t1) );
fim FAN_N1875_0 ( .fault(fault), .net(N1875), .FEN(FEN[1145]), .op(N1875_t0) );
fim FAN_N1875_1 ( .fault(fault), .net(N1875), .FEN(FEN[1146]), .op(N1875_t1) );
fim FAN_N2073_0 ( .fault(fault), .net(N2073), .FEN(FEN[1147]), .op(N2073_t0) );
fim FAN_N2073_1 ( .fault(fault), .net(N2073), .FEN(FEN[1148]), .op(N2073_t1) );
fim FAN_N3128_0 ( .fault(fault), .net(N3128), .FEN(FEN[1149]), .op(N3128_t0) );
fim FAN_N3128_1 ( .fault(fault), .net(N3128), .FEN(FEN[1150]), .op(N3128_t1) );
fim FAN_N3131_0 ( .fault(fault), .net(N3131), .FEN(FEN[1151]), .op(N3131_t0) );
fim FAN_N3131_1 ( .fault(fault), .net(N3131), .FEN(FEN[1152]), .op(N3131_t1) );
fim FAN_N3135_0 ( .fault(fault), .net(N3135), .FEN(FEN[1153]), .op(N3135_t0) );
fim FAN_N3135_1 ( .fault(fault), .net(N3135), .FEN(FEN[1154]), .op(N3135_t1) );
fim FAN_N3138_0 ( .fault(fault), .net(N3138), .FEN(FEN[1155]), .op(N3138_t0) );
fim FAN_N3138_1 ( .fault(fault), .net(N3138), .FEN(FEN[1156]), .op(N3138_t1) );
fim FAN_N3142_0 ( .fault(fault), .net(N3142), .FEN(FEN[1157]), .op(N3142_t0) );
fim FAN_N3142_1 ( .fault(fault), .net(N3142), .FEN(FEN[1158]), .op(N3142_t1) );
fim FAN_N3145_0 ( .fault(fault), .net(N3145), .FEN(FEN[1159]), .op(N3145_t0) );
fim FAN_N3145_1 ( .fault(fault), .net(N3145), .FEN(FEN[1160]), .op(N3145_t1) );
fim FAN_N3149_0 ( .fault(fault), .net(N3149), .FEN(FEN[1161]), .op(N3149_t0) );
fim FAN_N3149_1 ( .fault(fault), .net(N3149), .FEN(FEN[1162]), .op(N3149_t1) );
fim FAN_N1895_0 ( .fault(fault), .net(N1895), .FEN(FEN[1163]), .op(N1895_t0) );
fim FAN_N1895_1 ( .fault(fault), .net(N1895), .FEN(FEN[1164]), .op(N1895_t1) );
fim FAN_N2093_0 ( .fault(fault), .net(N2093), .FEN(FEN[1165]), .op(N2093_t0) );
fim FAN_N2093_1 ( .fault(fault), .net(N2093), .FEN(FEN[1166]), .op(N2093_t1) );
fim FAN_N3158_0 ( .fault(fault), .net(N3158), .FEN(FEN[1167]), .op(N3158_t0) );
fim FAN_N3158_1 ( .fault(fault), .net(N3158), .FEN(FEN[1168]), .op(N3158_t1) );
fim FAN_N3161_0 ( .fault(fault), .net(N3161), .FEN(FEN[1169]), .op(N3161_t0) );
fim FAN_N3161_1 ( .fault(fault), .net(N3161), .FEN(FEN[1170]), .op(N3161_t1) );
fim FAN_N3165_0 ( .fault(fault), .net(N3165), .FEN(FEN[1171]), .op(N3165_t0) );
fim FAN_N3165_1 ( .fault(fault), .net(N3165), .FEN(FEN[1172]), .op(N3165_t1) );
fim FAN_N3168_0 ( .fault(fault), .net(N3168), .FEN(FEN[1173]), .op(N3168_t0) );
fim FAN_N3168_1 ( .fault(fault), .net(N3168), .FEN(FEN[1174]), .op(N3168_t1) );
fim FAN_N2967_0 ( .fault(fault), .net(N2967), .FEN(FEN[1175]), .op(N2967_t0) );
fim FAN_N2967_1 ( .fault(fault), .net(N2967), .FEN(FEN[1176]), .op(N2967_t1) );
fim FAN_N2970_0 ( .fault(fault), .net(N2970), .FEN(FEN[1177]), .op(N2970_t0) );
fim FAN_N2970_1 ( .fault(fault), .net(N2970), .FEN(FEN[1178]), .op(N2970_t1) );
fim FAN_N3172_0 ( .fault(fault), .net(N3172), .FEN(FEN[1179]), .op(N3172_t0) );
fim FAN_N3172_1 ( .fault(fault), .net(N3172), .FEN(FEN[1180]), .op(N3172_t1) );
fim FAN_N3175_0 ( .fault(fault), .net(N3175), .FEN(FEN[1181]), .op(N3175_t0) );
fim FAN_N3175_1 ( .fault(fault), .net(N3175), .FEN(FEN[1182]), .op(N3175_t1) );
fim FAN_N3178_0 ( .fault(fault), .net(N3178), .FEN(FEN[1183]), .op(N3178_t0) );
fim FAN_N3178_1 ( .fault(fault), .net(N3178), .FEN(FEN[1184]), .op(N3178_t1) );
fim FAN_N3181_0 ( .fault(fault), .net(N3181), .FEN(FEN[1185]), .op(N3181_t0) );
fim FAN_N3181_1 ( .fault(fault), .net(N3181), .FEN(FEN[1186]), .op(N3181_t1) );
fim FAN_N3184_0 ( .fault(fault), .net(N3184), .FEN(FEN[1187]), .op(N3184_t0) );
fim FAN_N3184_1 ( .fault(fault), .net(N3184), .FEN(FEN[1188]), .op(N3184_t1) );
fim FAN_N3187_0 ( .fault(fault), .net(N3187), .FEN(FEN[1189]), .op(N3187_t0) );
fim FAN_N3187_1 ( .fault(fault), .net(N3187), .FEN(FEN[1190]), .op(N3187_t1) );
fim FAN_N3478_0 ( .fault(fault), .net(N3478), .FEN(FEN[1191]), .op(N3478_t0) );
fim FAN_N3478_1 ( .fault(fault), .net(N3478), .FEN(FEN[1192]), .op(N3478_t1) );
fim FAN_N3481_0 ( .fault(fault), .net(N3481), .FEN(FEN[1193]), .op(N3481_t0) );
fim FAN_N3481_1 ( .fault(fault), .net(N3481), .FEN(FEN[1194]), .op(N3481_t1) );
fim FAN_N3487_0 ( .fault(fault), .net(N3487), .FEN(FEN[1195]), .op(N3487_t0) );
fim FAN_N3487_1 ( .fault(fault), .net(N3487), .FEN(FEN[1196]), .op(N3487_t1) );
fim FAN_N3484_0 ( .fault(fault), .net(N3484), .FEN(FEN[1197]), .op(N3484_t0) );
fim FAN_N3484_1 ( .fault(fault), .net(N3484), .FEN(FEN[1198]), .op(N3484_t1) );
fim FAN_N3472_0 ( .fault(fault), .net(N3472), .FEN(FEN[1199]), .op(N3472_t0) );
fim FAN_N3472_1 ( .fault(fault), .net(N3472), .FEN(FEN[1200]), .op(N3472_t1) );
fim FAN_N3475_0 ( .fault(fault), .net(N3475), .FEN(FEN[1201]), .op(N3475_t0) );
fim FAN_N3475_1 ( .fault(fault), .net(N3475), .FEN(FEN[1202]), .op(N3475_t1) );
fim FAN_N3407_0 ( .fault(fault), .net(N3407), .FEN(FEN[1203]), .op(N3407_t0) );
fim FAN_N3407_1 ( .fault(fault), .net(N3407), .FEN(FEN[1204]), .op(N3407_t1) );
fim FAN_N3410_0 ( .fault(fault), .net(N3410), .FEN(FEN[1205]), .op(N3410_t0) );
fim FAN_N3410_1 ( .fault(fault), .net(N3410), .FEN(FEN[1206]), .op(N3410_t1) );
fim FAN_N3415_0 ( .fault(fault), .net(N3415), .FEN(FEN[1207]), .op(N3415_t0) );
fim FAN_N3415_1 ( .fault(fault), .net(N3415), .FEN(FEN[1208]), .op(N3415_t1) );
fim FAN_N3415_2 ( .fault(fault), .net(N3415), .FEN(FEN[1209]), .op(N3415_t2) );
fim FAN_N3122_0 ( .fault(fault), .net(N3122), .FEN(FEN[1210]), .op(N3122_t0) );
fim FAN_N3122_1 ( .fault(fault), .net(N3122), .FEN(FEN[1211]), .op(N3122_t1) );
fim FAN_N3125_0 ( .fault(fault), .net(N3125), .FEN(FEN[1212]), .op(N3125_t0) );
fim FAN_N3125_1 ( .fault(fault), .net(N3125), .FEN(FEN[1213]), .op(N3125_t1) );
fim FAN_N3419_0 ( .fault(fault), .net(N3419), .FEN(FEN[1214]), .op(N3419_t0) );
fim FAN_N3419_1 ( .fault(fault), .net(N3419), .FEN(FEN[1215]), .op(N3419_t1) );
fim FAN_N3419_2 ( .fault(fault), .net(N3419), .FEN(FEN[1216]), .op(N3419_t2) );
fim FAN_N3423_0 ( .fault(fault), .net(N3423), .FEN(FEN[1217]), .op(N3423_t0) );
fim FAN_N3423_1 ( .fault(fault), .net(N3423), .FEN(FEN[1218]), .op(N3423_t1) );
fim FAN_N3426_0 ( .fault(fault), .net(N3426), .FEN(FEN[1219]), .op(N3426_t0) );
fim FAN_N3426_1 ( .fault(fault), .net(N3426), .FEN(FEN[1220]), .op(N3426_t1) );
fim FAN_N3431_0 ( .fault(fault), .net(N3431), .FEN(FEN[1221]), .op(N3431_t0) );
fim FAN_N3431_1 ( .fault(fault), .net(N3431), .FEN(FEN[1222]), .op(N3431_t1) );
fim FAN_N3434_0 ( .fault(fault), .net(N3434), .FEN(FEN[1223]), .op(N3434_t0) );
fim FAN_N3434_1 ( .fault(fault), .net(N3434), .FEN(FEN[1224]), .op(N3434_t1) );
fim FAN_N3439_0 ( .fault(fault), .net(N3439), .FEN(FEN[1225]), .op(N3439_t0) );
fim FAN_N3439_1 ( .fault(fault), .net(N3439), .FEN(FEN[1226]), .op(N3439_t1) );
fim FAN_N3442_0 ( .fault(fault), .net(N3442), .FEN(FEN[1227]), .op(N3442_t0) );
fim FAN_N3442_1 ( .fault(fault), .net(N3442), .FEN(FEN[1228]), .op(N3442_t1) );
fim FAN_N3447_0 ( .fault(fault), .net(N3447), .FEN(FEN[1229]), .op(N3447_t0) );
fim FAN_N3447_1 ( .fault(fault), .net(N3447), .FEN(FEN[1230]), .op(N3447_t1) );
fim FAN_N3447_2 ( .fault(fault), .net(N3447), .FEN(FEN[1231]), .op(N3447_t2) );
fim FAN_N3152_0 ( .fault(fault), .net(N3152), .FEN(FEN[1232]), .op(N3152_t0) );
fim FAN_N3152_1 ( .fault(fault), .net(N3152), .FEN(FEN[1233]), .op(N3152_t1) );
fim FAN_N3155_0 ( .fault(fault), .net(N3155), .FEN(FEN[1234]), .op(N3155_t0) );
fim FAN_N3155_1 ( .fault(fault), .net(N3155), .FEN(FEN[1235]), .op(N3155_t1) );
fim FAN_N3451_0 ( .fault(fault), .net(N3451), .FEN(FEN[1236]), .op(N3451_t0) );
fim FAN_N3451_1 ( .fault(fault), .net(N3451), .FEN(FEN[1237]), .op(N3451_t1) );
fim FAN_N3451_2 ( .fault(fault), .net(N3451), .FEN(FEN[1238]), .op(N3451_t2) );
fim FAN_N3455_0 ( .fault(fault), .net(N3455), .FEN(FEN[1239]), .op(N3455_t0) );
fim FAN_N3455_1 ( .fault(fault), .net(N3455), .FEN(FEN[1240]), .op(N3455_t1) );
fim FAN_N3458_0 ( .fault(fault), .net(N3458), .FEN(FEN[1241]), .op(N3458_t0) );
fim FAN_N3458_1 ( .fault(fault), .net(N3458), .FEN(FEN[1242]), .op(N3458_t1) );
fim FAN_N3463_0 ( .fault(fault), .net(N3463), .FEN(FEN[1243]), .op(N3463_t0) );
fim FAN_N3463_1 ( .fault(fault), .net(N3463), .FEN(FEN[1244]), .op(N3463_t1) );
fim FAN_N3466_0 ( .fault(fault), .net(N3466), .FEN(FEN[1245]), .op(N3466_t0) );
fim FAN_N3466_1 ( .fault(fault), .net(N3466), .FEN(FEN[1246]), .op(N3466_t1) );
fim FAN_N3493_0 ( .fault(fault), .net(N3493), .FEN(FEN[1247]), .op(N3493_t0) );
fim FAN_N3493_1 ( .fault(fault), .net(N3493), .FEN(FEN[1248]), .op(N3493_t1) );
fim FAN_N3496_0 ( .fault(fault), .net(N3496), .FEN(FEN[1249]), .op(N3496_t0) );
fim FAN_N3496_1 ( .fault(fault), .net(N3496), .FEN(FEN[1250]), .op(N3496_t1) );
fim FAN_N3499_0 ( .fault(fault), .net(N3499), .FEN(FEN[1251]), .op(N3499_t0) );
fim FAN_N3499_1 ( .fault(fault), .net(N3499), .FEN(FEN[1252]), .op(N3499_t1) );
fim FAN_N3502_0 ( .fault(fault), .net(N3502), .FEN(FEN[1253]), .op(N3502_t0) );
fim FAN_N3502_1 ( .fault(fault), .net(N3502), .FEN(FEN[1254]), .op(N3502_t1) );
fim FAN_N3505_0 ( .fault(fault), .net(N3505), .FEN(FEN[1255]), .op(N3505_t0) );
fim FAN_N3505_1 ( .fault(fault), .net(N3505), .FEN(FEN[1256]), .op(N3505_t1) );
fim FAN_N3511_0 ( .fault(fault), .net(N3511), .FEN(FEN[1257]), .op(N3511_t0) );
fim FAN_N3511_1 ( .fault(fault), .net(N3511), .FEN(FEN[1258]), .op(N3511_t1) );
fim FAN_N3517_0 ( .fault(fault), .net(N3517), .FEN(FEN[1259]), .op(N3517_t0) );
fim FAN_N3517_1 ( .fault(fault), .net(N3517), .FEN(FEN[1260]), .op(N3517_t1) );
fim FAN_N3520_0 ( .fault(fault), .net(N3520), .FEN(FEN[1261]), .op(N3520_t0) );
fim FAN_N3520_1 ( .fault(fault), .net(N3520), .FEN(FEN[1262]), .op(N3520_t1) );
fim FAN_N3523_0 ( .fault(fault), .net(N3523), .FEN(FEN[1263]), .op(N3523_t0) );
fim FAN_N3523_1 ( .fault(fault), .net(N3523), .FEN(FEN[1264]), .op(N3523_t1) );
fim FAN_N3514_0 ( .fault(fault), .net(N3514), .FEN(FEN[1265]), .op(N3514_t0) );
fim FAN_N3514_1 ( .fault(fault), .net(N3514), .FEN(FEN[1266]), .op(N3514_t1) );
fim FAN_N3384_0 ( .fault(fault), .net(N3384), .FEN(FEN[1267]), .op(N3384_t0) );
fim FAN_N3384_1 ( .fault(fault), .net(N3384), .FEN(FEN[1268]), .op(N3384_t1) );
fim FAN_N3490_0 ( .fault(fault), .net(N3490), .FEN(FEN[1269]), .op(N3490_t0) );
fim FAN_N3490_1 ( .fault(fault), .net(N3490), .FEN(FEN[1270]), .op(N3490_t1) );
fim FAN_N3508_0 ( .fault(fault), .net(N3508), .FEN(FEN[1271]), .op(N3508_t0) );
fim FAN_N3508_1 ( .fault(fault), .net(N3508), .FEN(FEN[1272]), .op(N3508_t1) );
fim FAN_N3700_0 ( .fault(fault), .net(N3700), .FEN(FEN[1273]), .op(N3700_t0) );
fim FAN_N3700_1 ( .fault(fault), .net(N3700), .FEN(FEN[1274]), .op(N3700_t1) );
fim FAN_N3697_0 ( .fault(fault), .net(N3697), .FEN(FEN[1275]), .op(N3697_t0) );
fim FAN_N3697_1 ( .fault(fault), .net(N3697), .FEN(FEN[1276]), .op(N3697_t1) );
fim FAN_N3645_0 ( .fault(fault), .net(N3645), .FEN(FEN[1277]), .op(N3645_t0) );
fim FAN_N3645_1 ( .fault(fault), .net(N3645), .FEN(FEN[1278]), .op(N3645_t1) );
fim FAN_N3648_0 ( .fault(fault), .net(N3648), .FEN(FEN[1279]), .op(N3648_t0) );
fim FAN_N3648_1 ( .fault(fault), .net(N3648), .FEN(FEN[1280]), .op(N3648_t1) );
fim FAN_N3664_0 ( .fault(fault), .net(N3664), .FEN(FEN[1281]), .op(N3664_t0) );
fim FAN_N3664_1 ( .fault(fault), .net(N3664), .FEN(FEN[1282]), .op(N3664_t1) );
fim FAN_N3667_0 ( .fault(fault), .net(N3667), .FEN(FEN[1283]), .op(N3667_t0) );
fim FAN_N3667_1 ( .fault(fault), .net(N3667), .FEN(FEN[1284]), .op(N3667_t1) );
fim FAN_N3654_0 ( .fault(fault), .net(N3654), .FEN(FEN[1285]), .op(N3654_t0) );
fim FAN_N3654_1 ( .fault(fault), .net(N3654), .FEN(FEN[1286]), .op(N3654_t1) );
fim FAN_N3658_0 ( .fault(fault), .net(N3658), .FEN(FEN[1287]), .op(N3658_t0) );
fim FAN_N3658_1 ( .fault(fault), .net(N3658), .FEN(FEN[1288]), .op(N3658_t1) );
fim FAN_N3673_0 ( .fault(fault), .net(N3673), .FEN(FEN[1289]), .op(N3673_t0) );
fim FAN_N3673_1 ( .fault(fault), .net(N3673), .FEN(FEN[1290]), .op(N3673_t1) );
fim FAN_N1926_0 ( .fault(fault), .net(N1926), .FEN(FEN[1291]), .op(N1926_t0) );
fim FAN_N1926_1 ( .fault(fault), .net(N1926), .FEN(FEN[1292]), .op(N1926_t1) );
fim FAN_N1926_2 ( .fault(fault), .net(N1926), .FEN(FEN[1293]), .op(N1926_t2) );
fim FAN_N3677_0 ( .fault(fault), .net(N3677), .FEN(FEN[1294]), .op(N3677_t0) );
fim FAN_N3677_1 ( .fault(fault), .net(N3677), .FEN(FEN[1295]), .op(N3677_t1) );
fim FAN_N3682_0 ( .fault(fault), .net(N3682), .FEN(FEN[1296]), .op(N3682_t0) );
fim FAN_N3682_1 ( .fault(fault), .net(N3682), .FEN(FEN[1297]), .op(N3682_t1) );
fim FAN_N3690_0 ( .fault(fault), .net(N3690), .FEN(FEN[1298]), .op(N3690_t0) );
fim FAN_N3690_1 ( .fault(fault), .net(N3690), .FEN(FEN[1299]), .op(N3690_t1) );
fim FAN_N3721_0 ( .fault(fault), .net(N3721), .FEN(FEN[1300]), .op(N3721_t0) );
fim FAN_N3721_1 ( .fault(fault), .net(N3721), .FEN(FEN[1301]), .op(N3721_t1) );
fim FAN_N3721_2 ( .fault(fault), .net(N3721), .FEN(FEN[1302]), .op(N3721_t2) );
fim FAN_N3721_3 ( .fault(fault), .net(N3721), .FEN(FEN[1303]), .op(N3721_t3) );
fim FAN_N3721_4 ( .fault(fault), .net(N3721), .FEN(FEN[1304]), .op(N3721_t4) );
fim FAN_N3734_0 ( .fault(fault), .net(N3734), .FEN(FEN[1305]), .op(N3734_t0) );
fim FAN_N3734_1 ( .fault(fault), .net(N3734), .FEN(FEN[1306]), .op(N3734_t1) );
fim FAN_N3734_2 ( .fault(fault), .net(N3734), .FEN(FEN[1307]), .op(N3734_t2) );
fim FAN_N3740_0 ( .fault(fault), .net(N3740), .FEN(FEN[1308]), .op(N3740_t0) );
fim FAN_N3740_1 ( .fault(fault), .net(N3740), .FEN(FEN[1309]), .op(N3740_t1) );
fim FAN_N3743_0 ( .fault(fault), .net(N3743), .FEN(FEN[1310]), .op(N3743_t0) );
fim FAN_N3743_1 ( .fault(fault), .net(N3743), .FEN(FEN[1311]), .op(N3743_t1) );
fim FAN_N3743_2 ( .fault(fault), .net(N3743), .FEN(FEN[1312]), .op(N3743_t2) );
fim FAN_N3743_3 ( .fault(fault), .net(N3743), .FEN(FEN[1313]), .op(N3743_t3) );
fim FAN_N3743_4 ( .fault(fault), .net(N3743), .FEN(FEN[1314]), .op(N3743_t4) );
fim FAN_N3756_0 ( .fault(fault), .net(N3756), .FEN(FEN[1315]), .op(N3756_t0) );
fim FAN_N3756_1 ( .fault(fault), .net(N3756), .FEN(FEN[1316]), .op(N3756_t1) );
fim FAN_N3756_2 ( .fault(fault), .net(N3756), .FEN(FEN[1317]), .op(N3756_t2) );
fim FAN_N3762_0 ( .fault(fault), .net(N3762), .FEN(FEN[1318]), .op(N3762_t0) );
fim FAN_N3762_1 ( .fault(fault), .net(N3762), .FEN(FEN[1319]), .op(N3762_t1) );
fim FAN_N3786_0 ( .fault(fault), .net(N3786), .FEN(FEN[1320]), .op(N3786_t0) );
fim FAN_N3786_1 ( .fault(fault), .net(N3786), .FEN(FEN[1321]), .op(N3786_t1) );
fim FAN_N3800_0 ( .fault(fault), .net(N3800), .FEN(FEN[1322]), .op(N3800_t0) );
fim FAN_N3800_1 ( .fault(fault), .net(N3800), .FEN(FEN[1323]), .op(N3800_t1) );
fim FAN_N3821_0 ( .fault(fault), .net(N3821), .FEN(FEN[1324]), .op(N3821_t0) );
fim FAN_N3821_1 ( .fault(fault), .net(N3821), .FEN(FEN[1325]), .op(N3821_t1) );
fim FAN_N3824_0 ( .fault(fault), .net(N3824), .FEN(FEN[1326]), .op(N3824_t0) );
fim FAN_N3824_1 ( .fault(fault), .net(N3824), .FEN(FEN[1327]), .op(N3824_t1) );
fim FAN_N3830_0 ( .fault(fault), .net(N3830), .FEN(FEN[1328]), .op(N3830_t0) );
fim FAN_N3830_1 ( .fault(fault), .net(N3830), .FEN(FEN[1329]), .op(N3830_t1) );
fim FAN_N3827_0 ( .fault(fault), .net(N3827), .FEN(FEN[1330]), .op(N3827_t0) );
fim FAN_N3827_1 ( .fault(fault), .net(N3827), .FEN(FEN[1331]), .op(N3827_t1) );
fim FAN_N3812_0 ( .fault(fault), .net(N3812), .FEN(FEN[1332]), .op(N3812_t0) );
fim FAN_N3812_1 ( .fault(fault), .net(N3812), .FEN(FEN[1333]), .op(N3812_t1) );
fim FAN_N3818_0 ( .fault(fault), .net(N3818), .FEN(FEN[1334]), .op(N3818_t0) );
fim FAN_N3818_1 ( .fault(fault), .net(N3818), .FEN(FEN[1335]), .op(N3818_t1) );
fim FAN_N3809_0 ( .fault(fault), .net(N3809), .FEN(FEN[1336]), .op(N3809_t0) );
fim FAN_N3809_1 ( .fault(fault), .net(N3809), .FEN(FEN[1337]), .op(N3809_t1) );
fim FAN_N3838_0 ( .fault(fault), .net(N3838), .FEN(FEN[1338]), .op(N3838_t0) );
fim FAN_N3838_1 ( .fault(fault), .net(N3838), .FEN(FEN[1339]), .op(N3838_t1) );
fim FAN_N3838_2 ( .fault(fault), .net(N3838), .FEN(FEN[1340]), .op(N3838_t2) );
fim FAN_N3838_3 ( .fault(fault), .net(N3838), .FEN(FEN[1341]), .op(N3838_t3) );
fim FAN_N3845_0 ( .fault(fault), .net(N3845), .FEN(FEN[1342]), .op(N3845_t0) );
fim FAN_N3845_1 ( .fault(fault), .net(N3845), .FEN(FEN[1343]), .op(N3845_t1) );
fim FAN_N3845_2 ( .fault(fault), .net(N3845), .FEN(FEN[1344]), .op(N3845_t2) );
fim FAN_N3845_3 ( .fault(fault), .net(N3845), .FEN(FEN[1345]), .op(N3845_t3) );
fim FAN_N3850_0 ( .fault(fault), .net(N3850), .FEN(FEN[1346]), .op(N3850_t0) );
fim FAN_N3850_1 ( .fault(fault), .net(N3850), .FEN(FEN[1347]), .op(N3850_t1) );
fim FAN_N3855_0 ( .fault(fault), .net(N3855), .FEN(FEN[1348]), .op(N3855_t0) );
fim FAN_N3855_1 ( .fault(fault), .net(N3855), .FEN(FEN[1349]), .op(N3855_t1) );
fim FAN_N3858_0 ( .fault(fault), .net(N3858), .FEN(FEN[1350]), .op(N3858_t0) );
fim FAN_N3858_1 ( .fault(fault), .net(N3858), .FEN(FEN[1351]), .op(N3858_t1) );
fim FAN_N3861_0 ( .fault(fault), .net(N3861), .FEN(FEN[1352]), .op(N3861_t0) );
fim FAN_N3861_1 ( .fault(fault), .net(N3861), .FEN(FEN[1353]), .op(N3861_t1) );
fim FAN_N3865_0 ( .fault(fault), .net(N3865), .FEN(FEN[1354]), .op(N3865_t0) );
fim FAN_N3865_1 ( .fault(fault), .net(N3865), .FEN(FEN[1355]), .op(N3865_t1) );
fim FAN_N3868_0 ( .fault(fault), .net(N3868), .FEN(FEN[1356]), .op(N3868_t0) );
fim FAN_N3868_1 ( .fault(fault), .net(N3868), .FEN(FEN[1357]), .op(N3868_t1) );
fim FAN_N3921_0 ( .fault(fault), .net(N3921), .FEN(FEN[1358]), .op(N3921_t0) );
fim FAN_N3921_1 ( .fault(fault), .net(N3921), .FEN(FEN[1359]), .op(N3921_t1) );
fim FAN_N3932_0 ( .fault(fault), .net(N3932), .FEN(FEN[1360]), .op(N3932_t0) );
fim FAN_N3932_1 ( .fault(fault), .net(N3932), .FEN(FEN[1361]), .op(N3932_t1) );
fim FAN_N3926_0 ( .fault(fault), .net(N3926), .FEN(FEN[1362]), .op(N3926_t0) );
fim FAN_N3926_1 ( .fault(fault), .net(N3926), .FEN(FEN[1363]), .op(N3926_t1) );
fim FAN_N3926_2 ( .fault(fault), .net(N3926), .FEN(FEN[1364]), .op(N3926_t2) );
fim FAN_N3953_0 ( .fault(fault), .net(N3953), .FEN(FEN[1365]), .op(N3953_t0) );
fim FAN_N3953_1 ( .fault(fault), .net(N3953), .FEN(FEN[1366]), .op(N3953_t1) );
fim FAN_N3959_0 ( .fault(fault), .net(N3959), .FEN(FEN[1367]), .op(N3959_t0) );
fim FAN_N3959_1 ( .fault(fault), .net(N3959), .FEN(FEN[1368]), .op(N3959_t1) );
fim FAN_N3965_0 ( .fault(fault), .net(N3965), .FEN(FEN[1369]), .op(N3965_t0) );
fim FAN_N3965_1 ( .fault(fault), .net(N3965), .FEN(FEN[1370]), .op(N3965_t1) );
fim FAN_N3971_0 ( .fault(fault), .net(N3971), .FEN(FEN[1371]), .op(N3971_t0) );
fim FAN_N3971_1 ( .fault(fault), .net(N3971), .FEN(FEN[1372]), .op(N3971_t1) );
fim FAN_N3977_0 ( .fault(fault), .net(N3977), .FEN(FEN[1373]), .op(N3977_t0) );
fim FAN_N3977_1 ( .fault(fault), .net(N3977), .FEN(FEN[1374]), .op(N3977_t1) );
fim FAN_N3983_0 ( .fault(fault), .net(N3983), .FEN(FEN[1375]), .op(N3983_t0) );
fim FAN_N3983_1 ( .fault(fault), .net(N3983), .FEN(FEN[1376]), .op(N3983_t1) );
fim FAN_N3956_0 ( .fault(fault), .net(N3956), .FEN(FEN[1377]), .op(N3956_t0) );
fim FAN_N3956_1 ( .fault(fault), .net(N3956), .FEN(FEN[1378]), .op(N3956_t1) );
fim FAN_N3962_0 ( .fault(fault), .net(N3962), .FEN(FEN[1379]), .op(N3962_t0) );
fim FAN_N3962_1 ( .fault(fault), .net(N3962), .FEN(FEN[1380]), .op(N3962_t1) );
fim FAN_N3980_0 ( .fault(fault), .net(N3980), .FEN(FEN[1381]), .op(N3980_t0) );
fim FAN_N3980_1 ( .fault(fault), .net(N3980), .FEN(FEN[1382]), .op(N3980_t1) );
fim FAN_N3974_0 ( .fault(fault), .net(N3974), .FEN(FEN[1383]), .op(N3974_t0) );
fim FAN_N3974_1 ( .fault(fault), .net(N3974), .FEN(FEN[1384]), .op(N3974_t1) );
fim FAN_N3950_0 ( .fault(fault), .net(N3950), .FEN(FEN[1385]), .op(N3950_t0) );
fim FAN_N3950_1 ( .fault(fault), .net(N3950), .FEN(FEN[1386]), .op(N3950_t1) );
fim FAN_N3937_0 ( .fault(fault), .net(N3937), .FEN(FEN[1387]), .op(N3937_t0) );
fim FAN_N3937_1 ( .fault(fault), .net(N3937), .FEN(FEN[1388]), .op(N3937_t1) );
fim FAN_N3968_0 ( .fault(fault), .net(N3968), .FEN(FEN[1389]), .op(N3968_t0) );
fim FAN_N3968_1 ( .fault(fault), .net(N3968), .FEN(FEN[1390]), .op(N3968_t1) );
fim FAN_N3940_0 ( .fault(fault), .net(N3940), .FEN(FEN[1391]), .op(N3940_t0) );
fim FAN_N3940_1 ( .fault(fault), .net(N3940), .FEN(FEN[1392]), .op(N3940_t1) );
fim FAN_N3996_0 ( .fault(fault), .net(N3996), .FEN(FEN[1393]), .op(N3996_t0) );
fim FAN_N3996_1 ( .fault(fault), .net(N3996), .FEN(FEN[1394]), .op(N3996_t1) );
fim FAN_N3992_0 ( .fault(fault), .net(N3992), .FEN(FEN[1395]), .op(N3992_t0) );
fim FAN_N3992_1 ( .fault(fault), .net(N3992), .FEN(FEN[1396]), .op(N3992_t1) );
fim FAN_N4062_0 ( .fault(fault), .net(N4062), .FEN(FEN[1397]), .op(N4062_t0) );
fim FAN_N4062_1 ( .fault(fault), .net(N4062), .FEN(FEN[1398]), .op(N4062_t1) );
fim FAN_N4070_0 ( .fault(fault), .net(N4070), .FEN(FEN[1399]), .op(N4070_t0) );
fim FAN_N4070_1 ( .fault(fault), .net(N4070), .FEN(FEN[1400]), .op(N4070_t1) );
fim FAN_N4059_0 ( .fault(fault), .net(N4059), .FEN(FEN[1401]), .op(N4059_t0) );
fim FAN_N4059_1 ( .fault(fault), .net(N4059), .FEN(FEN[1402]), .op(N4059_t1) );
fim FAN_N4067_0 ( .fault(fault), .net(N4067), .FEN(FEN[1403]), .op(N4067_t0) );
fim FAN_N4067_1 ( .fault(fault), .net(N4067), .FEN(FEN[1404]), .op(N4067_t1) );
fim FAN_N4091_0 ( .fault(fault), .net(N4091), .FEN(FEN[1405]), .op(N4091_t0) );
fim FAN_N4091_1 ( .fault(fault), .net(N4091), .FEN(FEN[1406]), .op(N4091_t1) );
fim FAN_N4094_0 ( .fault(fault), .net(N4094), .FEN(FEN[1407]), .op(N4094_t0) );
fim FAN_N4094_1 ( .fault(fault), .net(N4094), .FEN(FEN[1408]), .op(N4094_t1) );
fim FAN_N4094_2 ( .fault(fault), .net(N4094), .FEN(FEN[1409]), .op(N4094_t2) );
fim FAN_N4116_0 ( .fault(fault), .net(N4116), .FEN(FEN[1410]), .op(N4116_t0) );
fim FAN_N4116_1 ( .fault(fault), .net(N4116), .FEN(FEN[1411]), .op(N4116_t1) );
fim FAN_N4119_0 ( .fault(fault), .net(N4119), .FEN(FEN[1412]), .op(N4119_t0) );
fim FAN_N4119_1 ( .fault(fault), .net(N4119), .FEN(FEN[1413]), .op(N4119_t1) );
fim FAN_N4123_0 ( .fault(fault), .net(N4123), .FEN(FEN[1414]), .op(N4123_t0) );
fim FAN_N4123_1 ( .fault(fault), .net(N4123), .FEN(FEN[1415]), .op(N4123_t1) );
fim FAN_N4128_0 ( .fault(fault), .net(N4128), .FEN(FEN[1416]), .op(N4128_t0) );
fim FAN_N4128_1 ( .fault(fault), .net(N4128), .FEN(FEN[1417]), .op(N4128_t1) );
fim FAN_N4128_2 ( .fault(fault), .net(N4128), .FEN(FEN[1418]), .op(N4128_t2) );
fim FAN_N4128_3 ( .fault(fault), .net(N4128), .FEN(FEN[1419]), .op(N4128_t3) );
fim FAN_N4128_4 ( .fault(fault), .net(N4128), .FEN(FEN[1420]), .op(N4128_t4) );
fim FAN_N3917_0 ( .fault(fault), .net(N3917), .FEN(FEN[1421]), .op(N3917_t0) );
fim FAN_N3917_1 ( .fault(fault), .net(N3917), .FEN(FEN[1422]), .op(N3917_t1) );
fim FAN_N4139_0 ( .fault(fault), .net(N4139), .FEN(FEN[1423]), .op(N4139_t0) );
fim FAN_N4139_1 ( .fault(fault), .net(N4139), .FEN(FEN[1424]), .op(N4139_t1) );
fim FAN_N4142_0 ( .fault(fault), .net(N4142), .FEN(FEN[1425]), .op(N4142_t0) );
fim FAN_N4142_1 ( .fault(fault), .net(N4142), .FEN(FEN[1426]), .op(N4142_t1) );
fim FAN_N4167_0 ( .fault(fault), .net(N4167), .FEN(FEN[1427]), .op(N4167_t0) );
fim FAN_N4167_1 ( .fault(fault), .net(N4167), .FEN(FEN[1428]), .op(N4167_t1) );
fim FAN_N4167_2 ( .fault(fault), .net(N4167), .FEN(FEN[1429]), .op(N4167_t2) );
fim FAN_N4167_3 ( .fault(fault), .net(N4167), .FEN(FEN[1430]), .op(N4167_t3) );
fim FAN_N4167_4 ( .fault(fault), .net(N4167), .FEN(FEN[1431]), .op(N4167_t4) );
fim FAN_N4167_5 ( .fault(fault), .net(N4167), .FEN(FEN[1432]), .op(N4167_t5) );
fim FAN_N4035_0 ( .fault(fault), .net(N4035), .FEN(FEN[1433]), .op(N4035_t0) );
fim FAN_N4035_1 ( .fault(fault), .net(N4035), .FEN(FEN[1434]), .op(N4035_t1) );
fim FAN_N4174_0 ( .fault(fault), .net(N4174), .FEN(FEN[1435]), .op(N4174_t0) );
fim FAN_N4174_1 ( .fault(fault), .net(N4174), .FEN(FEN[1436]), .op(N4174_t1) );
fim FAN_N4174_2 ( .fault(fault), .net(N4174), .FEN(FEN[1437]), .op(N4174_t2) );
fim FAN_N4174_3 ( .fault(fault), .net(N4174), .FEN(FEN[1438]), .op(N4174_t3) );
fim FAN_N3815_0 ( .fault(fault), .net(N3815), .FEN(FEN[1439]), .op(N3815_t0) );
fim FAN_N3815_1 ( .fault(fault), .net(N3815), .FEN(FEN[1440]), .op(N3815_t1) );
fim FAN_N4186_0 ( .fault(fault), .net(N4186), .FEN(FEN[1441]), .op(N4186_t0) );
fim FAN_N4186_1 ( .fault(fault), .net(N4186), .FEN(FEN[1442]), .op(N4186_t1) );
fim FAN_N4182_0 ( .fault(fault), .net(N4182), .FEN(FEN[1443]), .op(N4182_t0) );
fim FAN_N4182_1 ( .fault(fault), .net(N4182), .FEN(FEN[1444]), .op(N4182_t1) );
fim FAN_N4197_0 ( .fault(fault), .net(N4197), .FEN(FEN[1445]), .op(N4197_t0) );
fim FAN_N4197_1 ( .fault(fault), .net(N4197), .FEN(FEN[1446]), .op(N4197_t1) );
fim FAN_N4213_0 ( .fault(fault), .net(N4213), .FEN(FEN[1447]), .op(N4213_t0) );
fim FAN_N4213_1 ( .fault(fault), .net(N4213), .FEN(FEN[1448]), .op(N4213_t1) );
fim FAN_N4213_2 ( .fault(fault), .net(N4213), .FEN(FEN[1449]), .op(N4213_t2) );
fim FAN_N4213_3 ( .fault(fault), .net(N4213), .FEN(FEN[1450]), .op(N4213_t3) );
fim FAN_N4203_0 ( .fault(fault), .net(N4203), .FEN(FEN[1451]), .op(N4203_t0) );
fim FAN_N4203_1 ( .fault(fault), .net(N4203), .FEN(FEN[1452]), .op(N4203_t1) );
fim FAN_N4203_2 ( .fault(fault), .net(N4203), .FEN(FEN[1453]), .op(N4203_t2) );
fim FAN_N4203_3 ( .fault(fault), .net(N4203), .FEN(FEN[1454]), .op(N4203_t3) );
fim FAN_N4203_4 ( .fault(fault), .net(N4203), .FEN(FEN[1455]), .op(N4203_t4) );
fim FAN_N4209_0 ( .fault(fault), .net(N4209), .FEN(FEN[1456]), .op(N4209_t0) );
fim FAN_N4209_1 ( .fault(fault), .net(N4209), .FEN(FEN[1457]), .op(N4209_t1) );
fim FAN_N4209_2 ( .fault(fault), .net(N4209), .FEN(FEN[1458]), .op(N4209_t2) );
fim FAN_N4223_0 ( .fault(fault), .net(N4223), .FEN(FEN[1459]), .op(N4223_t0) );
fim FAN_N4223_1 ( .fault(fault), .net(N4223), .FEN(FEN[1460]), .op(N4223_t1) );
fim FAN_N4223_2 ( .fault(fault), .net(N4223), .FEN(FEN[1461]), .op(N4223_t2) );
fim FAN_N4223_3 ( .fault(fault), .net(N4223), .FEN(FEN[1462]), .op(N4223_t3) );
fim FAN_N4218_0 ( .fault(fault), .net(N4218), .FEN(FEN[1463]), .op(N4218_t0) );
fim FAN_N4218_1 ( .fault(fault), .net(N4218), .FEN(FEN[1464]), .op(N4218_t1) );
fim FAN_N4218_2 ( .fault(fault), .net(N4218), .FEN(FEN[1465]), .op(N4218_t2) );
fim FAN_N4218_3 ( .fault(fault), .net(N4218), .FEN(FEN[1466]), .op(N4218_t3) );
fim FAN_N3913_0 ( .fault(fault), .net(N3913), .FEN(FEN[1467]), .op(N3913_t0) );
fim FAN_N3913_1 ( .fault(fault), .net(N3913), .FEN(FEN[1468]), .op(N3913_t1) );
fim FAN_N4247_0 ( .fault(fault), .net(N4247), .FEN(FEN[1469]), .op(N4247_t0) );
fim FAN_N4247_1 ( .fault(fault), .net(N4247), .FEN(FEN[1470]), .op(N4247_t1) );
fim FAN_N4242_0 ( .fault(fault), .net(N4242), .FEN(FEN[1471]), .op(N4242_t0) );
fim FAN_N4242_1 ( .fault(fault), .net(N4242), .FEN(FEN[1472]), .op(N4242_t1) );
fim FAN_N4287_0 ( .fault(fault), .net(N4287), .FEN(FEN[1473]), .op(N4287_t0) );
fim FAN_N4287_1 ( .fault(fault), .net(N4287), .FEN(FEN[1474]), .op(N4287_t1) );
fim FAN_N4287_2 ( .fault(fault), .net(N4287), .FEN(FEN[1475]), .op(N4287_t2) );
fim FAN_N4284_0 ( .fault(fault), .net(N4284), .FEN(FEN[1476]), .op(N4284_t0) );
fim FAN_N4284_1 ( .fault(fault), .net(N4284), .FEN(FEN[1477]), .op(N4284_t1) );
fim FAN_N4331_0 ( .fault(fault), .net(N4331), .FEN(FEN[1478]), .op(N4331_t0) );
fim FAN_N4331_1 ( .fault(fault), .net(N4331), .FEN(FEN[1479]), .op(N4331_t1) );
fim FAN_N4296_0 ( .fault(fault), .net(N4296), .FEN(FEN[1480]), .op(N4296_t0) );
fim FAN_N4296_1 ( .fault(fault), .net(N4296), .FEN(FEN[1481]), .op(N4296_t1) );
fim FAN_N4305_0 ( .fault(fault), .net(N4305), .FEN(FEN[1482]), .op(N4305_t0) );
fim FAN_N4305_1 ( .fault(fault), .net(N4305), .FEN(FEN[1483]), .op(N4305_t1) );
fim FAN_N4305_2 ( .fault(fault), .net(N4305), .FEN(FEN[1484]), .op(N4305_t2) );
fim FAN_N4305_3 ( .fault(fault), .net(N4305), .FEN(FEN[1485]), .op(N4305_t3) );
fim FAN_N4200_0 ( .fault(fault), .net(N4200), .FEN(FEN[1486]), .op(N4200_t0) );
fim FAN_N4200_1 ( .fault(fault), .net(N4200), .FEN(FEN[1487]), .op(N4200_t1) );
fim FAN_N4356_0 ( .fault(fault), .net(N4356), .FEN(FEN[1488]), .op(N4356_t0) );
fim FAN_N4356_1 ( .fault(fault), .net(N4356), .FEN(FEN[1489]), .op(N4356_t1) );
fim FAN_N4365_0 ( .fault(fault), .net(N4365), .FEN(FEN[1490]), .op(N4365_t0) );
fim FAN_N4365_1 ( .fault(fault), .net(N4365), .FEN(FEN[1491]), .op(N4365_t1) );
fim FAN_N4368_0 ( .fault(fault), .net(N4368), .FEN(FEN[1492]), .op(N4368_t0) );
fim FAN_N4368_1 ( .fault(fault), .net(N4368), .FEN(FEN[1493]), .op(N4368_t1) );
fim FAN_N4371_0 ( .fault(fault), .net(N4371), .FEN(FEN[1494]), .op(N4371_t0) );
fim FAN_N4371_1 ( .fault(fault), .net(N4371), .FEN(FEN[1495]), .op(N4371_t1) );
fim FAN_N4310_0 ( .fault(fault), .net(N4310), .FEN(FEN[1496]), .op(N4310_t0) );
fim FAN_N4310_1 ( .fault(fault), .net(N4310), .FEN(FEN[1497]), .op(N4310_t1) );
fim FAN_N4310_2 ( .fault(fault), .net(N4310), .FEN(FEN[1498]), .op(N4310_t2) );
fim FAN_N4353_0 ( .fault(fault), .net(N4353), .FEN(FEN[1499]), .op(N4353_t0) );
fim FAN_N4353_1 ( .fault(fault), .net(N4353), .FEN(FEN[1500]), .op(N4353_t1) );
fim FAN_N4359_0 ( .fault(fault), .net(N4359), .FEN(FEN[1501]), .op(N4359_t0) );
fim FAN_N4359_1 ( .fault(fault), .net(N4359), .FEN(FEN[1502]), .op(N4359_t1) );
fim FAN_N4362_0 ( .fault(fault), .net(N4362), .FEN(FEN[1503]), .op(N4362_t0) );
fim FAN_N4362_1 ( .fault(fault), .net(N4362), .FEN(FEN[1504]), .op(N4362_t1) );
fim FAN_N4319_0 ( .fault(fault), .net(N4319), .FEN(FEN[1505]), .op(N4319_t0) );
fim FAN_N4319_1 ( .fault(fault), .net(N4319), .FEN(FEN[1506]), .op(N4319_t1) );
fim FAN_N4398_0 ( .fault(fault), .net(N4398), .FEN(FEN[1507]), .op(N4398_t0) );
fim FAN_N4398_1 ( .fault(fault), .net(N4398), .FEN(FEN[1508]), .op(N4398_t1) );
fim FAN_N4413_0 ( .fault(fault), .net(N4413), .FEN(FEN[1509]), .op(N4413_t0) );
fim FAN_N4413_1 ( .fault(fault), .net(N4413), .FEN(FEN[1510]), .op(N4413_t1) );
fim FAN_N4435_0 ( .fault(fault), .net(N4435), .FEN(FEN[1511]), .op(N4435_t0) );
fim FAN_N4435_1 ( .fault(fault), .net(N4435), .FEN(FEN[1512]), .op(N4435_t1) );
fim FAN_N4421_0 ( .fault(fault), .net(N4421), .FEN(FEN[1513]), .op(N4421_t0) );
fim FAN_N4421_1 ( .fault(fault), .net(N4421), .FEN(FEN[1514]), .op(N4421_t1) );
fim FAN_N4427_0 ( .fault(fault), .net(N4427), .FEN(FEN[1515]), .op(N4427_t0) );
fim FAN_N4427_1 ( .fault(fault), .net(N4427), .FEN(FEN[1516]), .op(N4427_t1) );
fim FAN_N4416_0 ( .fault(fault), .net(N4416), .FEN(FEN[1517]), .op(N4416_t0) );
fim FAN_N4416_1 ( .fault(fault), .net(N4416), .FEN(FEN[1518]), .op(N4416_t1) );
fim FAN_N4430_0 ( .fault(fault), .net(N4430), .FEN(FEN[1519]), .op(N4430_t0) );
fim FAN_N4430_1 ( .fault(fault), .net(N4430), .FEN(FEN[1520]), .op(N4430_t1) );
fim FAN_N4387_0 ( .fault(fault), .net(N4387), .FEN(FEN[1521]), .op(N4387_t0) );
fim FAN_N4387_1 ( .fault(fault), .net(N4387), .FEN(FEN[1522]), .op(N4387_t1) );
fim FAN_N4390_0 ( .fault(fault), .net(N4390), .FEN(FEN[1523]), .op(N4390_t0) );
fim FAN_N4390_1 ( .fault(fault), .net(N4390), .FEN(FEN[1524]), .op(N4390_t1) );
fim FAN_N4443_0 ( .fault(fault), .net(N4443), .FEN(FEN[1525]), .op(N4443_t0) );
fim FAN_N4443_1 ( .fault(fault), .net(N4443), .FEN(FEN[1526]), .op(N4443_t1) );
fim FAN_N4493_0 ( .fault(fault), .net(N4493), .FEN(FEN[1527]), .op(N4493_t0) );
fim FAN_N4493_1 ( .fault(fault), .net(N4493), .FEN(FEN[1528]), .op(N4493_t1) );
fim FAN_N4465_0 ( .fault(fault), .net(N4465), .FEN(FEN[1529]), .op(N4465_t0) );
fim FAN_N4465_1 ( .fault(fault), .net(N4465), .FEN(FEN[1530]), .op(N4465_t1) );
fim FAN_N4468_0 ( .fault(fault), .net(N4468), .FEN(FEN[1531]), .op(N4468_t0) );
fim FAN_N4468_1 ( .fault(fault), .net(N4468), .FEN(FEN[1532]), .op(N4468_t1) );
fim FAN_N4479_0 ( .fault(fault), .net(N4479), .FEN(FEN[1533]), .op(N4479_t0) );
fim FAN_N4479_1 ( .fault(fault), .net(N4479), .FEN(FEN[1534]), .op(N4479_t1) );
fim FAN_N4458_0 ( .fault(fault), .net(N4458), .FEN(FEN[1535]), .op(N4458_t0) );
fim FAN_N4458_1 ( .fault(fault), .net(N4458), .FEN(FEN[1536]), .op(N4458_t1) );
fim FAN_N2758_0 ( .fault(fault), .net(N2758), .FEN(FEN[1537]), .op(N2758_t0) );
fim FAN_N2758_1 ( .fault(fault), .net(N2758), .FEN(FEN[1538]), .op(N2758_t1) );
fim FAN_N4498_0 ( .fault(fault), .net(N4498), .FEN(FEN[1539]), .op(N4498_t0) );
fim FAN_N4498_1 ( .fault(fault), .net(N4498), .FEN(FEN[1540]), .op(N4498_t1) );
fim FAN_N2761_0 ( .fault(fault), .net(N2761), .FEN(FEN[1541]), .op(N2761_t0) );
fim FAN_N2761_1 ( .fault(fault), .net(N2761), .FEN(FEN[1542]), .op(N2761_t1) );
fim FAN_N4531_0 ( .fault(fault), .net(N4531), .FEN(FEN[1543]), .op(N4531_t0) );
fim FAN_N4531_1 ( .fault(fault), .net(N4531), .FEN(FEN[1544]), .op(N4531_t1) );
fim FAN_N4534_0 ( .fault(fault), .net(N4534), .FEN(FEN[1545]), .op(N4534_t0) );
fim FAN_N4534_1 ( .fault(fault), .net(N4534), .FEN(FEN[1546]), .op(N4534_t1) );
fim FAN_N4537_0 ( .fault(fault), .net(N4537), .FEN(FEN[1547]), .op(N4537_t0) );
fim FAN_N4537_1 ( .fault(fault), .net(N4537), .FEN(FEN[1548]), .op(N4537_t1) );
fim FAN_N4540_0 ( .fault(fault), .net(N4540), .FEN(FEN[1549]), .op(N4540_t0) );
fim FAN_N4540_1 ( .fault(fault), .net(N4540), .FEN(FEN[1550]), .op(N4540_t1) );
fim FAN_N4503_0 ( .fault(fault), .net(N4503), .FEN(FEN[1551]), .op(N4503_t0) );
fim FAN_N4503_1 ( .fault(fault), .net(N4503), .FEN(FEN[1552]), .op(N4503_t1) );
fim FAN_N4569_0 ( .fault(fault), .net(N4569), .FEN(FEN[1553]), .op(N4569_t0) );
fim FAN_N4569_1 ( .fault(fault), .net(N4569), .FEN(FEN[1554]), .op(N4569_t1) );
fim FAN_N4576_0 ( .fault(fault), .net(N4576), .FEN(FEN[1555]), .op(N4576_t0) );
fim FAN_N4576_1 ( .fault(fault), .net(N4576), .FEN(FEN[1556]), .op(N4576_t1) );
fim FAN_N4581_0 ( .fault(fault), .net(N4581), .FEN(FEN[1557]), .op(N4581_t0) );
fim FAN_N4581_1 ( .fault(fault), .net(N4581), .FEN(FEN[1558]), .op(N4581_t1) );
fim FAN_N4584_0 ( .fault(fault), .net(N4584), .FEN(FEN[1559]), .op(N4584_t0) );
fim FAN_N4584_1 ( .fault(fault), .net(N4584), .FEN(FEN[1560]), .op(N4584_t1) );
fim FAN_N4559_0 ( .fault(fault), .net(N4559), .FEN(FEN[1561]), .op(N4559_t0) );
fim FAN_N4559_1 ( .fault(fault), .net(N4559), .FEN(FEN[1562]), .op(N4559_t1) );
fim FAN_N4549_0 ( .fault(fault), .net(N4549), .FEN(FEN[1563]), .op(N4549_t0) );
fim FAN_N4549_1 ( .fault(fault), .net(N4549), .FEN(FEN[1564]), .op(N4549_t1) );
fim FAN_N4564_0 ( .fault(fault), .net(N4564), .FEN(FEN[1565]), .op(N4564_t0) );
fim FAN_N4564_1 ( .fault(fault), .net(N4564), .FEN(FEN[1566]), .op(N4564_t1) );
fim FAN_N4564_2 ( .fault(fault), .net(N4564), .FEN(FEN[1567]), .op(N4564_t2) );
fim FAN_N4616_0 ( .fault(fault), .net(N4616), .FEN(FEN[1568]), .op(N4616_t0) );
fim FAN_N4616_1 ( .fault(fault), .net(N4616), .FEN(FEN[1569]), .op(N4616_t1) );
fim FAN_N4619_0 ( .fault(fault), .net(N4619), .FEN(FEN[1570]), .op(N4619_t0) );
fim FAN_N4619_1 ( .fault(fault), .net(N4619), .FEN(FEN[1571]), .op(N4619_t1) );
fim FAN_N4623_0 ( .fault(fault), .net(N4623), .FEN(FEN[1572]), .op(N4623_t0) );
fim FAN_N4623_1 ( .fault(fault), .net(N4623), .FEN(FEN[1573]), .op(N4623_t1) );
fim FAN_N4613_0 ( .fault(fault), .net(N4613), .FEN(FEN[1574]), .op(N4613_t0) );
fim FAN_N4613_1 ( .fault(fault), .net(N4613), .FEN(FEN[1575]), .op(N4613_t1) );
fim FAN_N4593_0 ( .fault(fault), .net(N4593), .FEN(FEN[1576]), .op(N4593_t0) );
fim FAN_N4593_1 ( .fault(fault), .net(N4593), .FEN(FEN[1577]), .op(N4593_t1) );
fim FAN_N4599_0 ( .fault(fault), .net(N4599), .FEN(FEN[1578]), .op(N4599_t0) );
fim FAN_N4599_1 ( .fault(fault), .net(N4599), .FEN(FEN[1579]), .op(N4599_t1) );
fim FAN_N4656_0 ( .fault(fault), .net(N4656), .FEN(FEN[1580]), .op(N4656_t0) );
fim FAN_N4656_1 ( .fault(fault), .net(N4656), .FEN(FEN[1581]), .op(N4656_t1) );
fim FAN_N4659_0 ( .fault(fault), .net(N4659), .FEN(FEN[1582]), .op(N4659_t0) );
fim FAN_N4659_1 ( .fault(fault), .net(N4659), .FEN(FEN[1583]), .op(N4659_t1) );
fim FAN_N4644_0 ( .fault(fault), .net(N4644), .FEN(FEN[1584]), .op(N4644_t0) );
fim FAN_N4644_1 ( .fault(fault), .net(N4644), .FEN(FEN[1585]), .op(N4644_t1) );
fim FAN_N4664_0 ( .fault(fault), .net(N4664), .FEN(FEN[1586]), .op(N4664_t0) );
fim FAN_N4664_1 ( .fault(fault), .net(N4664), .FEN(FEN[1587]), .op(N4664_t1) );
fim FAN_N4647_0 ( .fault(fault), .net(N4647), .FEN(FEN[1588]), .op(N4647_t0) );
fim FAN_N4647_1 ( .fault(fault), .net(N4647), .FEN(FEN[1589]), .op(N4647_t1) );
fim FAN_N4650_0 ( .fault(fault), .net(N4650), .FEN(FEN[1590]), .op(N4650_t0) );
fim FAN_N4650_1 ( .fault(fault), .net(N4650), .FEN(FEN[1591]), .op(N4650_t1) );
fim FAN_N4350_0 ( .fault(fault), .net(N4350), .FEN(FEN[1592]), .op(N4350_t0) );
fim FAN_N4350_1 ( .fault(fault), .net(N4350), .FEN(FEN[1593]), .op(N4350_t1) );
fim FAN_N4691_0 ( .fault(fault), .net(N4691), .FEN(FEN[1594]), .op(N4691_t0) );
fim FAN_N4691_1 ( .fault(fault), .net(N4691), .FEN(FEN[1595]), .op(N4691_t1) );
fim FAN_N4694_0 ( .fault(fault), .net(N4694), .FEN(FEN[1596]), .op(N4694_t0) );
fim FAN_N4694_1 ( .fault(fault), .net(N4694), .FEN(FEN[1597]), .op(N4694_t1) );
fim FAN_N4697_0 ( .fault(fault), .net(N4697), .FEN(FEN[1598]), .op(N4697_t0) );
fim FAN_N4697_1 ( .fault(fault), .net(N4697), .FEN(FEN[1599]), .op(N4697_t1) );
fim FAN_N4700_0 ( .fault(fault), .net(N4700), .FEN(FEN[1600]), .op(N4700_t0) );
fim FAN_N4700_1 ( .fault(fault), .net(N4700), .FEN(FEN[1601]), .op(N4700_t1) );
fim FAN_N4730_0 ( .fault(fault), .net(N4730), .FEN(FEN[1602]), .op(N4730_t0) );
fim FAN_N4730_1 ( .fault(fault), .net(N4730), .FEN(FEN[1603]), .op(N4730_t1) );
fim FAN_N4711_0 ( .fault(fault), .net(N4711), .FEN(FEN[1604]), .op(N4711_t0) );
fim FAN_N4711_1 ( .fault(fault), .net(N4711), .FEN(FEN[1605]), .op(N4711_t1) );
fim FAN_N4717_0 ( .fault(fault), .net(N4717), .FEN(FEN[1606]), .op(N4717_t0) );
fim FAN_N4717_1 ( .fault(fault), .net(N4717), .FEN(FEN[1607]), .op(N4717_t1) );
fim FAN_N4717_2 ( .fault(fault), .net(N4717), .FEN(FEN[1608]), .op(N4717_t2) );
fim FAN_N4722_0 ( .fault(fault), .net(N4722), .FEN(FEN[1609]), .op(N4722_t0) );
fim FAN_N4722_1 ( .fault(fault), .net(N4722), .FEN(FEN[1610]), .op(N4722_t1) );
fim FAN_N4722_2 ( .fault(fault), .net(N4722), .FEN(FEN[1611]), .op(N4722_t2) );
fim FAN_N4727_0 ( .fault(fault), .net(N4727), .FEN(FEN[1612]), .op(N4727_t0) );
fim FAN_N4727_1 ( .fault(fault), .net(N4727), .FEN(FEN[1613]), .op(N4727_t1) );
fim FAN_N4769_0 ( .fault(fault), .net(N4769), .FEN(FEN[1614]), .op(N4769_t0) );
fim FAN_N4769_1 ( .fault(fault), .net(N4769), .FEN(FEN[1615]), .op(N4769_t1) );
fim FAN_N4772_0 ( .fault(fault), .net(N4772), .FEN(FEN[1616]), .op(N4772_t0) );
fim FAN_N4772_1 ( .fault(fault), .net(N4772), .FEN(FEN[1617]), .op(N4772_t1) );
fim FAN_N4775_0 ( .fault(fault), .net(N4775), .FEN(FEN[1618]), .op(N4775_t0) );
fim FAN_N4775_1 ( .fault(fault), .net(N4775), .FEN(FEN[1619]), .op(N4775_t1) );
fim FAN_N4743_0 ( .fault(fault), .net(N4743), .FEN(FEN[1620]), .op(N4743_t0) );
fim FAN_N4743_1 ( .fault(fault), .net(N4743), .FEN(FEN[1621]), .op(N4743_t1) );
fim FAN_N4743_2 ( .fault(fault), .net(N4743), .FEN(FEN[1622]), .op(N4743_t2) );
fim FAN_N4757_0 ( .fault(fault), .net(N4757), .FEN(FEN[1623]), .op(N4757_t0) );
fim FAN_N4757_1 ( .fault(fault), .net(N4757), .FEN(FEN[1624]), .op(N4757_t1) );
fim FAN_N4757_2 ( .fault(fault), .net(N4757), .FEN(FEN[1625]), .op(N4757_t2) );
fim FAN_N4740_0 ( .fault(fault), .net(N4740), .FEN(FEN[1626]), .op(N4740_t0) );
fim FAN_N4740_1 ( .fault(fault), .net(N4740), .FEN(FEN[1627]), .op(N4740_t1) );
fim FAN_N4805_0 ( .fault(fault), .net(N4805), .FEN(FEN[1628]), .op(N4805_t0) );
fim FAN_N4805_1 ( .fault(fault), .net(N4805), .FEN(FEN[1629]), .op(N4805_t1) );
fim FAN_N4808_0 ( .fault(fault), .net(N4808), .FEN(FEN[1630]), .op(N4808_t0) );
fim FAN_N4808_1 ( .fault(fault), .net(N4808), .FEN(FEN[1631]), .op(N4808_t1) );
fim FAN_N4794_0 ( .fault(fault), .net(N4794), .FEN(FEN[1632]), .op(N4794_t0) );
fim FAN_N4794_1 ( .fault(fault), .net(N4794), .FEN(FEN[1633]), .op(N4794_t1) );
fim FAN_N4797_0 ( .fault(fault), .net(N4797), .FEN(FEN[1634]), .op(N4797_t0) );
fim FAN_N4797_1 ( .fault(fault), .net(N4797), .FEN(FEN[1635]), .op(N4797_t1) );
fim FAN_N4341_0 ( .fault(fault), .net(N4341), .FEN(FEN[1636]), .op(N4341_t0) );
fim FAN_N4341_1 ( .fault(fault), .net(N4341), .FEN(FEN[1637]), .op(N4341_t1) );
fim FAN_N4812_0 ( .fault(fault), .net(N4812), .FEN(FEN[1638]), .op(N4812_t0) );
fim FAN_N4812_1 ( .fault(fault), .net(N4812), .FEN(FEN[1639]), .op(N4812_t1) );
fim FAN_N4844_0 ( .fault(fault), .net(N4844), .FEN(FEN[1640]), .op(N4844_t0) );
fim FAN_N4844_1 ( .fault(fault), .net(N4844), .FEN(FEN[1641]), .op(N4844_t1) );
fim FAN_N4847_0 ( .fault(fault), .net(N4847), .FEN(FEN[1642]), .op(N4847_t0) );
fim FAN_N4847_1 ( .fault(fault), .net(N4847), .FEN(FEN[1643]), .op(N4847_t1) );
fim FAN_N4823_0 ( .fault(fault), .net(N4823), .FEN(FEN[1644]), .op(N4823_t0) );
fim FAN_N4823_1 ( .fault(fault), .net(N4823), .FEN(FEN[1645]), .op(N4823_t1) );
fim FAN_N4850_0 ( .fault(fault), .net(N4850), .FEN(FEN[1646]), .op(N4850_t0) );
fim FAN_N4850_1 ( .fault(fault), .net(N4850), .FEN(FEN[1647]), .op(N4850_t1) );
fim FAN_N4854_0 ( .fault(fault), .net(N4854), .FEN(FEN[1648]), .op(N4854_t0) );
fim FAN_N4854_1 ( .fault(fault), .net(N4854), .FEN(FEN[1649]), .op(N4854_t1) );
fim FAN_N4818_0 ( .fault(fault), .net(N4818), .FEN(FEN[1650]), .op(N4818_t0) );
fim FAN_N4818_1 ( .fault(fault), .net(N4818), .FEN(FEN[1651]), .op(N4818_t1) );
fim FAN_N4818_2 ( .fault(fault), .net(N4818), .FEN(FEN[1652]), .op(N4818_t2) );
fim FAN_N4880_0 ( .fault(fault), .net(N4880), .FEN(FEN[1653]), .op(N4880_t0) );
fim FAN_N4880_1 ( .fault(fault), .net(N4880), .FEN(FEN[1654]), .op(N4880_t1) );
fim FAN_N4889_0 ( .fault(fault), .net(N4889), .FEN(FEN[1655]), .op(N4889_t0) );
fim FAN_N4889_1 ( .fault(fault), .net(N4889), .FEN(FEN[1656]), .op(N4889_t1) );
fim FAN_N4876_0 ( .fault(fault), .net(N4876), .FEN(FEN[1657]), .op(N4876_t0) );
fim FAN_N4876_1 ( .fault(fault), .net(N4876), .FEN(FEN[1658]), .op(N4876_t1) );
fim FAN_N4876_2 ( .fault(fault), .net(N4876), .FEN(FEN[1659]), .op(N4876_t2) );
fim FAN_N4916_0 ( .fault(fault), .net(N4916), .FEN(FEN[1660]), .op(N4916_t0) );
fim FAN_N4916_1 ( .fault(fault), .net(N4916), .FEN(FEN[1661]), .op(N4916_t1) );
fim FAN_N2764_0 ( .fault(fault), .net(N2764), .FEN(FEN[1662]), .op(N2764_t0) );
fim FAN_N2764_1 ( .fault(fault), .net(N2764), .FEN(FEN[1663]), .op(N2764_t1) );
fim FAN_N2483_0 ( .fault(fault), .net(N2483), .FEN(FEN[1664]), .op(N2483_t0) );
fim FAN_N2483_1 ( .fault(fault), .net(N2483), .FEN(FEN[1665]), .op(N2483_t1) );
fim FAN_N4921_0 ( .fault(fault), .net(N4921), .FEN(FEN[1666]), .op(N4921_t0) );
fim FAN_N4921_1 ( .fault(fault), .net(N4921), .FEN(FEN[1667]), .op(N4921_t1) );
fim FAN_N4937_0 ( .fault(fault), .net(N4937), .FEN(FEN[1668]), .op(N4937_t0) );
fim FAN_N4937_1 ( .fault(fault), .net(N4937), .FEN(FEN[1669]), .op(N4937_t1) );
fim FAN_N4940_0 ( .fault(fault), .net(N4940), .FEN(FEN[1670]), .op(N4940_t0) );
fim FAN_N4940_1 ( .fault(fault), .net(N4940), .FEN(FEN[1671]), .op(N4940_t1) );
fim FAN_N4946_0 ( .fault(fault), .net(N4946), .FEN(FEN[1672]), .op(N4946_t0) );
fim FAN_N4946_1 ( .fault(fault), .net(N4946), .FEN(FEN[1673]), .op(N4946_t1) );
fim FAN_N4913_0 ( .fault(fault), .net(N4913), .FEN(FEN[1674]), .op(N4913_t0) );
fim FAN_N4913_1 ( .fault(fault), .net(N4913), .FEN(FEN[1675]), .op(N4913_t1) );
fim FAN_N4954_0 ( .fault(fault), .net(N4954), .FEN(FEN[1676]), .op(N4954_t0) );
fim FAN_N4954_1 ( .fault(fault), .net(N4954), .FEN(FEN[1677]), .op(N4954_t1) );
fim FAN_N4344_0 ( .fault(fault), .net(N4344), .FEN(FEN[1678]), .op(N4344_t0) );
fim FAN_N4344_1 ( .fault(fault), .net(N4344), .FEN(FEN[1679]), .op(N4344_t1) );
fim FAN_N4800_0 ( .fault(fault), .net(N4800), .FEN(FEN[1680]), .op(N4800_t0) );
fim FAN_N4800_1 ( .fault(fault), .net(N4800), .FEN(FEN[1681]), .op(N4800_t1) );
fim FAN_N4957_0 ( .fault(fault), .net(N4957), .FEN(FEN[1682]), .op(N4957_t0) );
fim FAN_N4957_1 ( .fault(fault), .net(N4957), .FEN(FEN[1683]), .op(N4957_t1) );
fim FAN_N4347_0 ( .fault(fault), .net(N4347), .FEN(FEN[1684]), .op(N4347_t0) );
fim FAN_N4347_1 ( .fault(fault), .net(N4347), .FEN(FEN[1685]), .op(N4347_t1) );
fim FAN_N4838_0 ( .fault(fault), .net(N4838), .FEN(FEN[1686]), .op(N4838_t0) );
fim FAN_N4838_1 ( .fault(fault), .net(N4838), .FEN(FEN[1687]), .op(N4838_t1) );
fim FAN_N4973_0 ( .fault(fault), .net(N4973), .FEN(FEN[1688]), .op(N4973_t0) );
fim FAN_N4973_1 ( .fault(fault), .net(N4973), .FEN(FEN[1689]), .op(N4973_t1) );
fim FAN_N4475_0 ( .fault(fault), .net(N4475), .FEN(FEN[1690]), .op(N4475_t0) );
fim FAN_N4475_1 ( .fault(fault), .net(N4475), .FEN(FEN[1691]), .op(N4475_t1) );
fim FAN_N4991_0 ( .fault(fault), .net(N4991), .FEN(FEN[1692]), .op(N4991_t0) );
fim FAN_N4991_1 ( .fault(fault), .net(N4991), .FEN(FEN[1693]), .op(N4991_t1) );
fim FAN_N4999_0 ( .fault(fault), .net(N4999), .FEN(FEN[1694]), .op(N4999_t0) );
fim FAN_N4999_1 ( .fault(fault), .net(N4999), .FEN(FEN[1695]), .op(N4999_t1) );
fim FAN_N4996_0 ( .fault(fault), .net(N4996), .FEN(FEN[1696]), .op(N4996_t0) );
fim FAN_N4996_1 ( .fault(fault), .net(N4996), .FEN(FEN[1697]), .op(N4996_t1) );
fim FAN_N4988_0 ( .fault(fault), .net(N4988), .FEN(FEN[1698]), .op(N4988_t0) );
fim FAN_N4988_1 ( .fault(fault), .net(N4988), .FEN(FEN[1699]), .op(N4988_t1) );
fim FAN_N5021_0 ( .fault(fault), .net(N5021), .FEN(FEN[1700]), .op(N5021_t0) );
fim FAN_N5021_1 ( .fault(fault), .net(N5021), .FEN(FEN[1701]), .op(N5021_t1) );
fim FAN_N4831_0 ( .fault(fault), .net(N4831), .FEN(FEN[1702]), .op(N4831_t0) );
fim FAN_N4831_1 ( .fault(fault), .net(N4831), .FEN(FEN[1703]), .op(N4831_t1) );
fim FAN_N5010_0 ( .fault(fault), .net(N5010), .FEN(FEN[1704]), .op(N5010_t0) );
fim FAN_N5010_1 ( .fault(fault), .net(N5010), .FEN(FEN[1705]), .op(N5010_t1) );
fim FAN_N4472_0 ( .fault(fault), .net(N4472), .FEN(FEN[1706]), .op(N4472_t0) );
fim FAN_N4472_1 ( .fault(fault), .net(N4472), .FEN(FEN[1707]), .op(N4472_t1) );
fim FAN_N4907_0 ( .fault(fault), .net(N4907), .FEN(FEN[1708]), .op(N4907_t0) );
fim FAN_N4907_1 ( .fault(fault), .net(N4907), .FEN(FEN[1709]), .op(N4907_t1) );
fim FAN_N5013_0 ( .fault(fault), .net(N5013), .FEN(FEN[1710]), .op(N5013_t0) );
fim FAN_N5013_1 ( .fault(fault), .net(N5013), .FEN(FEN[1711]), .op(N5013_t1) );
fim FAN_N4338_0 ( .fault(fault), .net(N4338), .FEN(FEN[1712]), .op(N4338_t0) );
fim FAN_N4338_1 ( .fault(fault), .net(N4338), .FEN(FEN[1713]), .op(N4338_t1) );
fim FAN_N5018_0 ( .fault(fault), .net(N5018), .FEN(FEN[1714]), .op(N5018_t0) );
fim FAN_N5018_1 ( .fault(fault), .net(N5018), .FEN(FEN[1715]), .op(N5018_t1) );
fim FAN_N4985_0 ( .fault(fault), .net(N4985), .FEN(FEN[1716]), .op(N4985_t0) );
fim FAN_N4985_1 ( .fault(fault), .net(N4985), .FEN(FEN[1717]), .op(N4985_t1) );
fim FAN_N5030_0 ( .fault(fault), .net(N5030), .FEN(FEN[1718]), .op(N5030_t0) );
fim FAN_N5030_1 ( .fault(fault), .net(N5030), .FEN(FEN[1719]), .op(N5030_t1) );
fim FAN_N4335_0 ( .fault(fault), .net(N4335), .FEN(FEN[1720]), .op(N4335_t0) );
fim FAN_N4335_1 ( .fault(fault), .net(N4335), .FEN(FEN[1721]), .op(N4335_t1) );
fim FAN_N5039_0 ( .fault(fault), .net(N5039), .FEN(FEN[1722]), .op(N5039_t0) );
fim FAN_N5039_1 ( .fault(fault), .net(N5039), .FEN(FEN[1723]), .op(N5039_t1) );
fim FAN_N5042_0 ( .fault(fault), .net(N5042), .FEN(FEN[1724]), .op(N5042_t0) );
fim FAN_N5042_1 ( .fault(fault), .net(N5042), .FEN(FEN[1725]), .op(N5042_t1) );
fim FAN_N5050_0 ( .fault(fault), .net(N5050), .FEN(FEN[1726]), .op(N5050_t0) );
fim FAN_N5050_1 ( .fault(fault), .net(N5050), .FEN(FEN[1727]), .op(N5050_t1) );
fim FAN_N5050_2 ( .fault(fault), .net(N5050), .FEN(FEN[1728]), .op(N5050_t2) );
fim FAN_N5050_3 ( .fault(fault), .net(N5050), .FEN(FEN[1729]), .op(N5050_t3) );
fim FAN_N5061_0 ( .fault(fault), .net(N5061), .FEN(FEN[1730]), .op(N5061_t0) );
fim FAN_N5061_1 ( .fault(fault), .net(N5061), .FEN(FEN[1731]), .op(N5061_t1) );
fim FAN_N5070_0 ( .fault(fault), .net(N5070), .FEN(FEN[1732]), .op(N5070_t0) );
fim FAN_N5070_1 ( .fault(fault), .net(N5070), .FEN(FEN[1733]), .op(N5070_t1) );
fim FAN_N5058_0 ( .fault(fault), .net(N5058), .FEN(FEN[1734]), .op(N5058_t0) );
fim FAN_N5058_1 ( .fault(fault), .net(N5058), .FEN(FEN[1735]), .op(N5058_t1) );
fim FAN_N1461_0 ( .fault(fault), .net(N1461), .FEN(FEN[1736]), .op(N1461_t0) );
fim FAN_N1461_1 ( .fault(fault), .net(N1461), .FEN(FEN[1737]), .op(N1461_t1) );
fim FAN_N5080_0 ( .fault(fault), .net(N5080), .FEN(FEN[1738]), .op(N5080_t0) );
fim FAN_N5080_1 ( .fault(fault), .net(N5080), .FEN(FEN[1739]), .op(N5080_t1) );
fim FAN_N5080_2 ( .fault(fault), .net(N5080), .FEN(FEN[1740]), .op(N5080_t2) );
fim FAN_N5080_3 ( .fault(fault), .net(N5080), .FEN(FEN[1741]), .op(N5080_t3) );
fim FAN_N5055_0 ( .fault(fault), .net(N5055), .FEN(FEN[1742]), .op(N5055_t0) );
fim FAN_N5055_1 ( .fault(fault), .net(N5055), .FEN(FEN[1743]), .op(N5055_t1) );
fim FAN_N5085_0 ( .fault(fault), .net(N5085), .FEN(FEN[1744]), .op(N5085_t0) );
fim FAN_N5085_1 ( .fault(fault), .net(N5085), .FEN(FEN[1745]), .op(N5085_t1) );
fim FAN_N5111_0 ( .fault(fault), .net(N5111), .FEN(FEN[1746]), .op(N5111_t0) );
fim FAN_N5111_1 ( .fault(fault), .net(N5111), .FEN(FEN[1747]), .op(N5111_t1) );
fim FAN_N5117_0 ( .fault(fault), .net(N5117), .FEN(FEN[1748]), .op(N5117_t0) );
fim FAN_N5117_1 ( .fault(fault), .net(N5117), .FEN(FEN[1749]), .op(N5117_t1) );
fim FAN_N5114_0 ( .fault(fault), .net(N5114), .FEN(FEN[1750]), .op(N5114_t0) );
fim FAN_N5114_1 ( .fault(fault), .net(N5114), .FEN(FEN[1751]), .op(N5114_t1) );
fim FAN_N5066_0 ( .fault(fault), .net(N5066), .FEN(FEN[1752]), .op(N5066_t0) );
fim FAN_N5066_1 ( .fault(fault), .net(N5066), .FEN(FEN[1753]), .op(N5066_t1) );
fim FAN_N5133_0 ( .fault(fault), .net(N5133), .FEN(FEN[1754]), .op(N5133_t0) );
fim FAN_N5133_1 ( .fault(fault), .net(N5133), .FEN(FEN[1755]), .op(N5133_t1) );
fim FAN_N5122_0 ( .fault(fault), .net(N5122), .FEN(FEN[1756]), .op(N5122_t0) );
fim FAN_N5122_1 ( .fault(fault), .net(N5122), .FEN(FEN[1757]), .op(N5122_t1) );
fim FAN_N5139_0 ( .fault(fault), .net(N5139), .FEN(FEN[1758]), .op(N5139_t0) );
fim FAN_N5139_1 ( .fault(fault), .net(N5139), .FEN(FEN[1759]), .op(N5139_t1) );
fim FAN_N5128_0 ( .fault(fault), .net(N5128), .FEN(FEN[1760]), .op(N5128_t0) );
fim FAN_N5128_1 ( .fault(fault), .net(N5128), .FEN(FEN[1761]), .op(N5128_t1) );
fim FAN_N5151_0 ( .fault(fault), .net(N5151), .FEN(FEN[1762]), .op(N5151_t0) );
fim FAN_N5151_1 ( .fault(fault), .net(N5151), .FEN(FEN[1763]), .op(N5151_t1) );
fim FAN_N5154_0 ( .fault(fault), .net(N5154), .FEN(FEN[1764]), .op(N5154_t0) );
fim FAN_N5154_1 ( .fault(fault), .net(N5154), .FEN(FEN[1765]), .op(N5154_t1) );
fim FAN_N5160_0 ( .fault(fault), .net(N5160), .FEN(FEN[1766]), .op(N5160_t0) );
fim FAN_N5160_1 ( .fault(fault), .net(N5160), .FEN(FEN[1767]), .op(N5160_t1) );
fim FAN_N5163_0 ( .fault(fault), .net(N5163), .FEN(FEN[1768]), .op(N5163_t0) );
fim FAN_N5163_1 ( .fault(fault), .net(N5163), .FEN(FEN[1769]), .op(N5163_t1) );
fim FAN_N5145_0 ( .fault(fault), .net(N5145), .FEN(FEN[1770]), .op(N5145_t0) );
fim FAN_N5145_1 ( .fault(fault), .net(N5145), .FEN(FEN[1771]), .op(N5145_t1) );
fim FAN_N5174_0 ( .fault(fault), .net(N5174), .FEN(FEN[1772]), .op(N5174_t0) );
fim FAN_N5174_1 ( .fault(fault), .net(N5174), .FEN(FEN[1773]), .op(N5174_t1) );
fim FAN_N5177_0 ( .fault(fault), .net(N5177), .FEN(FEN[1774]), .op(N5177_t0) );
fim FAN_N5177_1 ( .fault(fault), .net(N5177), .FEN(FEN[1775]), .op(N5177_t1) );
fim FAN_N5184_0 ( .fault(fault), .net(N5184), .FEN(FEN[1776]), .op(N5184_t0) );
fim FAN_N5184_1 ( .fault(fault), .net(N5184), .FEN(FEN[1777]), .op(N5184_t1) );
fim FAN_N5188_0 ( .fault(fault), .net(N5188), .FEN(FEN[1778]), .op(N5188_t0) );
fim FAN_N5188_1 ( .fault(fault), .net(N5188), .FEN(FEN[1779]), .op(N5188_t1) );
fim FAN_N5205_0 ( .fault(fault), .net(N5205), .FEN(FEN[1780]), .op(N5205_t0) );
fim FAN_N5205_1 ( .fault(fault), .net(N5205), .FEN(FEN[1781]), .op(N5205_t1) );
fim FAN_N5209_0 ( .fault(fault), .net(N5209), .FEN(FEN[1782]), .op(N5209_t0) );
fim FAN_N5209_1 ( .fault(fault), .net(N5209), .FEN(FEN[1783]), .op(N5209_t1) );
fim FAN_N5228_0 ( .fault(fault), .net(N5228), .FEN(FEN[1784]), .op(N5228_t0) );
fim FAN_N5228_1 ( .fault(fault), .net(N5228), .FEN(FEN[1785]), .op(N5228_t1) );
fim FAN_N5236_0 ( .fault(fault), .net(N5236), .FEN(FEN[1786]), .op(N5236_t0) );
fim FAN_N5236_1 ( .fault(fault), .net(N5236), .FEN(FEN[1787]), .op(N5236_t1) );
fim FAN_N5236_2 ( .fault(fault), .net(N5236), .FEN(FEN[1788]), .op(N5236_t2) );
fim FAN_N5254_0 ( .fault(fault), .net(N5254), .FEN(FEN[1789]), .op(N5254_t0) );
fim FAN_N5254_1 ( .fault(fault), .net(N5254), .FEN(FEN[1790]), .op(N5254_t1) );
fim FAN_N2307_0 ( .fault(fault), .net(N2307), .FEN(FEN[1791]), .op(N2307_t0) );
fim FAN_N2307_1 ( .fault(fault), .net(N2307), .FEN(FEN[1792]), .op(N2307_t1) );
fim FAN_N5250_0 ( .fault(fault), .net(N5250), .FEN(FEN[1793]), .op(N5250_t0) );
fim FAN_N5250_1 ( .fault(fault), .net(N5250), .FEN(FEN[1794]), .op(N5250_t1) );
fim FAN_N2310_0 ( .fault(fault), .net(N2310), .FEN(FEN[1795]), .op(N2310_t0) );
fim FAN_N2310_1 ( .fault(fault), .net(N2310), .FEN(FEN[1796]), .op(N2310_t1) );
fim FAN_N5269_0 ( .fault(fault), .net(N5269), .FEN(FEN[1797]), .op(N5269_t0) );
fim FAN_N5269_1 ( .fault(fault), .net(N5269), .FEN(FEN[1798]), .op(N5269_t1) );
fim FAN_N5266_0 ( .fault(fault), .net(N5266), .FEN(FEN[1799]), .op(N5266_t0) );
fim FAN_N5266_1 ( .fault(fault), .net(N5266), .FEN(FEN[1800]), .op(N5266_t1) );
fim FAN_N5258_0 ( .fault(fault), .net(N5258), .FEN(FEN[1801]), .op(N5258_t0) );
fim FAN_N5258_1 ( .fault(fault), .net(N5258), .FEN(FEN[1802]), .op(N5258_t1) );
fim FAN_N5279_0 ( .fault(fault), .net(N5279), .FEN(FEN[1803]), .op(N5279_t0) );
fim FAN_N5279_1 ( .fault(fault), .net(N5279), .FEN(FEN[1804]), .op(N5279_t1) );
fim FAN_N5292_0 ( .fault(fault), .net(N5292), .FEN(FEN[1805]), .op(N5292_t0) );
fim FAN_N5292_1 ( .fault(fault), .net(N5292), .FEN(FEN[1806]), .op(N5292_t1) );
fim FAN_N5289_0 ( .fault(fault), .net(N5289), .FEN(FEN[1807]), .op(N5289_t0) );
fim FAN_N5289_1 ( .fault(fault), .net(N5289), .FEN(FEN[1808]), .op(N5289_t1) );
fim FAN_N5306_0 ( .fault(fault), .net(N5306), .FEN(FEN[1809]), .op(N5306_t0) );
fim FAN_N5306_1 ( .fault(fault), .net(N5306), .FEN(FEN[1810]), .op(N5306_t1) );
fim FAN_N5303_0 ( .fault(fault), .net(N5303), .FEN(FEN[1811]), .op(N5303_t0) );
fim FAN_N5303_1 ( .fault(fault), .net(N5303), .FEN(FEN[1812]), .op(N5303_t1) );
fim FAN_N5298_0 ( .fault(fault), .net(N5298), .FEN(FEN[1813]), .op(N5298_t0) );
fim FAN_N5298_1 ( .fault(fault), .net(N5298), .FEN(FEN[1814]), .op(N5298_t1) );
fim FAN_N5309_0 ( .fault(fault), .net(N5309), .FEN(FEN[1815]), .op(N5309_t0) );
fim FAN_N5309_1 ( .fault(fault), .net(N5309), .FEN(FEN[1816]), .op(N5309_t1) );
fim FAN_N5324_0 ( .fault(fault), .net(N5324), .FEN(FEN[1817]), .op(N5324_t0) );
fim FAN_N5324_1 ( .fault(fault), .net(N5324), .FEN(FEN[1818]), .op(N5324_t1) );
fim FAN_N5327_0 ( .fault(fault), .net(N5327), .FEN(FEN[1819]), .op(N5327_t0) );
fim FAN_N5327_1 ( .fault(fault), .net(N5327), .FEN(FEN[1820]), .op(N5327_t1) );
fim FAN_N5332_0 ( .fault(fault), .net(N5332), .FEN(FEN[1821]), .op(N5332_t0) );
fim FAN_N5332_1 ( .fault(fault), .net(N5332), .FEN(FEN[1822]), .op(N5332_t1) );
fim FAN_N5335_0 ( .fault(fault), .net(N5335), .FEN(FEN[1823]), .op(N5335_t0) );
fim FAN_N5335_1 ( .fault(fault), .net(N5335), .FEN(FEN[1824]), .op(N5335_t1) );
initial begin
    FEN <= {1824'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {1824'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,1824'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,1824'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN <= {FEN[1823:0], FEN[1824]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
// EndFaultModel

//Anchor
buf BUFF1_1 (N655, N50_t0);
not NOT1_2 (N665, N50_t1);
buf BUFF1_3 (N670, N58_t0);
not NOT1_4 (N679, N58_t1);
buf BUFF1_5 (N683, N68_t0);
not NOT1_6 (N686, N68_t1);
buf BUFF1_7 (N690, N68_t2);
buf BUFF1_8 (N699, N77_t0);
not NOT1_9 (N702, N77_t1);
buf BUFF1_10 (N706, N77_t2);
buf BUFF1_11 (N715, N87_t0);
not NOT1_12 (N724, N87_t1);
buf BUFF1_13 (N727, N97_t0);
not NOT1_14 (N736, N97_t1);
buf BUFF1_15 (N740, N107_t0);
not NOT1_16 (N749, N107_t1);
buf BUFF1_17 (N753, N116_t0);
not NOT1_18 (N763, N116_t1);
or OR2_19 (N768, N257_t0, N264_t0);
not NOT1_20 (N769, N1_t0);
buf BUFF1_21 (N772, N1_t1);
not NOT1_22 (N779, N1_t2);
buf BUFF1_23 (N782, N13_t0);
not NOT1_24 (N786, N13_t1);
and AND2_25 (N793, N13_t2, N20_t0);
not NOT1_26 (N794, N20_t1);
buf BUFF1_27 (N798, N20_t2);
not NOT1_28 (N803, N20_t3);
not NOT1_29 (N820, N33_t0);
buf BUFF1_30 (N821, N33_t1);
not NOT1_31 (N825, N33_t2);
and AND2_32 (N829, N33_t3, N41_t0);
not NOT1_33 (N832, N41_t1);
or OR2_34 (N835, N41_t2, N45_t0);
buf BUFF1_35 (N836, N45_t1);
not NOT1_36 (N839, N45_t2);
not NOT1_37 (N842, N50_t2);
buf BUFF1_38 (N845, N58_t2);
not NOT1_39 (N848, N58_t3);
buf BUFF1_40 (N851, N68_t3);
not NOT1_41 (N854, N68_t4);
buf BUFF1_42 (N858, N87_t2);
not NOT1_43 (N861, N87_t3);
buf BUFF1_44 (N864, N97_t2);
not NOT1_45 (N867, N97_t3);
not NOT1_46 (N870, N107_t2);
buf BUFF1_47 (N874, N1_t3);
buf BUFF1_48 (N877, N68_t5);
buf BUFF1_49 (N880, N107_t3);
not NOT1_50 (N883, N20_t4);
buf BUFF1_51 (N886, N190_t0);
not NOT1_52 (N889, N200_t0);
and AND2_53 (N890, N20_t5, N200_t1);
nand NAND2_54 (N891, N20_t6, N200_t2);
and AND2_55 (N892, N20_t7, N179_t0);
not NOT1_56 (N895, N20_t8);
or OR2_57 (N896, N349_t, N33_t4);
nand NAND2_58 (N913, N1_t4, N13_t3);
nand NAND3_59 (N914, N1_t5, N20_t9, N33_t5);
not NOT1_60 (N915, N20_t10);
not NOT1_61 (N916, N33_t6);
buf BUFF1_62 (N917, N179_t1);
not NOT1_63 (N920, N213_t0);
buf BUFF1_64 (N923, N343_t0);
buf BUFF1_65 (N926, N226_t0);
buf BUFF1_66 (N929, N232_t0);
buf BUFF1_67 (N932, N238_t0);
buf BUFF1_68 (N935, N244_t0);
buf BUFF1_69 (N938, N250_t0);
buf BUFF1_70 (N941, N257_t1);
buf BUFF1_71 (N944, N264_t1);
buf BUFF1_72 (N947, N270_t0);
buf BUFF1_73 (N950, N50_t3);
buf BUFF1_74 (N953, N58_t4);
buf BUFF1_75 (N956, N58_t5);
buf BUFF1_76 (N959, N97_t4);
buf BUFF1_77 (N962, N97_t5);
buf BUFF1_78 (N965, N330_t0);
and AND2_79 (N1067, N250_t1, N768);
or OR2_80 (N1117, N820, N20_t11);
or OR2_81 (N1179, N895, N169_t0);
not NOT1_82 (N1196, N793);
or OR2_83 (N1197, N915, N1_t6);
and AND2_84 (N1202, N913, N914);
or OR2_85 (N1219, N916, N1_t7);
and AND3_86 (N1250, N842_t0, N848_t0, N854_t0);
nand NAND2_87 (N1251, N226_t1, N655_t0);
nand NAND2_88 (N1252, N232_t1, N670_t0);
nand NAND2_89 (N1253, N238_t1, N690_t0);
nand NAND2_90 (N1254, N244_t1, N706_t0);
nand NAND2_91 (N1255, N250_t2, N715_t0);
nand NAND2_92 (N1256, N257_t2, N727_t0);
nand NAND2_93 (N1257, N264_t2, N740_t0);
nand NAND2_94 (N1258, N270_t1, N753_t0);
not NOT1_95 (N1259, N926_t0);
not NOT1_96 (N1260, N929_t0);
not NOT1_97 (N1261, N932_t0);
not NOT1_98 (N1262, N935_t0);
nand NAND2_99 (N1263, N679_t0, N686_t0);
nand NAND2_100 (N1264, N736_t0, N749_t0);
nand NAND2_101 (N1267, N683_t0, N699_t0);
buf BUFF1_102 (N1268, N665_t0);
not NOT1_103 (N1271, N953_t0);
not NOT1_104 (N1272, N959_t0);
buf BUFF1_105 (N1273, N839_t0);
buf BUFF1_106 (N1276, N839_t1);
buf BUFF1_107 (N1279, N782_t0);
buf BUFF1_108 (N1298, N825_t0);
buf BUFF1_109 (N1302, N832_t0);
and AND2_110 (N1306, N779_t0, N835);
and AND3_111 (N1315, N779_t1, N836_t0, N832_t1);
and AND2_112 (N1322, N769_t0, N836_t1);
and AND3_113 (N1325, N772_t0, N786_t0, N798_t0);
nand NAND3_114 (N1328, N772_t1, N786_t1, N798_t1);
nand NAND2_115 (N1331, N772_t2, N786_t2);
buf BUFF1_116 (N1334, N874_t0);
nand NAND3_117 (N1337, N782_t1, N794_t0, N45_t3);
nand NAND3_118 (N1338, N842_t1, N848_t1, N854_t1);
not NOT1_119 (N1339, N956_t0);
and AND3_120 (N1340, N861_t0, N867_t0, N870_t0);
nand NAND3_121 (N1343, N861_t1, N867_t1, N870_t1);
not NOT1_122 (N1344, N962_t0);
not NOT1_123 (N1345, N803_t0);
not NOT1_124 (N1346, N803_t1);
not NOT1_125 (N1347, N803_t2);
not NOT1_126 (N1348, N803_t3);
not NOT1_127 (N1349, N803_t4);
not NOT1_128 (N1350, N803_t5);
not NOT1_129 (N1351, N803_t6);
not NOT1_130 (N1352, N803_t7);
or OR2_131 (N1353, N883_t0, N886_t0);
nor NOR2_132 (N1358, N883_t1, N886_t1);
buf BUFF1_133 (N1363, N892_t0);
not NOT1_134 (N1366, N892_t1);
buf BUFF1_135 (N1369, N821_t0);
buf BUFF1_136 (N1384, N825_t1);
not NOT1_137 (N1401, N896_t0);
not NOT1_138 (N1402, N896_t1);
not NOT1_139 (N1403, N896_t2);
not NOT1_140 (N1404, N896_t3);
not NOT1_141 (N1405, N896_t4);
not NOT1_142 (N1406, N896_t5);
not NOT1_143 (N1407, N896_t6);
not NOT1_144 (N1408, N896_t7);
or OR2_145 (N1409, N1_t8, N1196);
not NOT1_146 (N1426, N829_t0);
not NOT1_147 (N1427, N829_t1);
and AND3_148 (N1452, N769_t1, N782_t2, N794_t1);
not NOT1_149 (N1459, N917_t0);
not NOT1_150 (N1460, N965_t0);
or OR2_151 (N1461, N920_t0, N923_t0);
nor NOR2_152 (N1464, N920_t1, N923_t1);
not NOT1_153 (N1467, N938_t0);
not NOT1_154 (N1468, N941_t0);
not NOT1_155 (N1469, N944_t0);
not NOT1_156 (N1470, N947_t0);
buf BUFF1_157 (N1471, N679_t1);
not NOT1_158 (N1474, N950_t0);
buf BUFF1_159 (N1475, N686_t1);
buf BUFF1_160 (N1478, N702_t0);
buf BUFF1_161 (N1481, N724_t0);
buf BUFF1_162 (N1484, N736_t1);
buf BUFF1_163 (N1487, N749_t1);
buf BUFF1_164 (N1490, N763_t0);
buf BUFF1_165 (N1493, N877_t0);
buf BUFF1_166 (N1496, N877_t1);
buf BUFF1_167 (N1499, N880_t0);
buf BUFF1_168 (N1502, N880_t1);
nand NAND2_169 (N1505, N702_t1, N1250);
and AND4_170 (N1507, N1251, N1252, N1253, N1254);
and AND4_171 (N1508, N1255, N1256, N1257, N1258);
nand NAND2_172 (N1509, N929_t1, N1259);
nand NAND2_173 (N1510, N926_t1, N1260);
nand NAND2_174 (N1511, N935_t1, N1261);
nand NAND2_175 (N1512, N932_t1, N1262);
and AND2_176 (N1520, N655_t1, N1263);
and AND2_177 (N1562, N874_t1, N1337);
not NOT1_178 (N1579, N1117_t0);
and AND2_179 (N1580, N803_t8, N1117_t1);
and AND2_180 (N1581, N1338, N1345);
not NOT1_181 (N1582, N1117_t2);
and AND2_182 (N1583, N803_t9, N1117_t3);
not NOT1_183 (N1584, N1117_t4);
and AND2_184 (N1585, N803_t10, N1117_t5);
and AND2_185 (N1586, N854_t2, N1347);
not NOT1_186 (N1587, N1117_t6);
and AND2_187 (N1588, N803_t11, N1117_t7);
and AND2_188 (N1589, N77_t3, N1348);
not NOT1_189 (N1590, N1117_t8);
and AND2_190 (N1591, N803_t12, N1117_t9);
and AND2_191 (N1592, N1343, N1349);
not NOT1_192 (N1593, N1117_t10);
and AND2_193 (N1594, N803_t13, N1117_t11);
not NOT1_194 (N1595, N1117_t12);
and AND2_195 (N1596, N803_t14, N1117_t13);
and AND2_196 (N1597, N870_t2, N1351);
not NOT1_197 (N1598, N1117_t14);
and AND2_198 (N1599, N803_t15, N1117_t15);
and AND2_199 (N1600, N116_t2, N1352);
and AND2_200 (N1643, N222_t, N1401);
and AND2_201 (N1644, N223_t0, N1402);
and AND2_202 (N1645, N226_t2, N1403);
and AND2_203 (N1646, N232_t2, N1404);
and AND2_204 (N1647, N238_t2, N1405);
and AND2_205 (N1648, N244_t2, N1406);
and AND2_206 (N1649, N250_t3, N1407);
and AND2_207 (N1650, N257_t3, N1408);
and AND3_208 (N1667, N1_t9, N13_t4, N1426);
and AND3_209 (N1670, N1_t10, N13_t5, N1427);
not NOT1_210 (N1673, N1202_t0);
not NOT1_211 (N1674, N1202_t1);
not NOT1_212 (N1675, N1202_t2);
not NOT1_213 (N1676, N1202_t3);
not NOT1_214 (N1677, N1202_t4);
not NOT1_215 (N1678, N1202_t5);
not NOT1_216 (N1679, N1202_t6);
not NOT1_217 (N1680, N1202_t7);
nand NAND2_218 (N1691, N941_t1, N1467);
nand NAND2_219 (N1692, N938_t1, N1468);
nand NAND2_220 (N1693, N947_t1, N1469);
nand NAND2_221 (N1694, N944_t1, N1470);
not NOT1_222 (N1713, N1505);
and AND2_223 (N1714, N87_t4, N1264_t0);
nand NAND2_224 (N1715, N1509, N1510);
nand NAND2_225 (N1718, N1511, N1512);
nand NAND2_226 (N1721, N1507, N1508);
and AND2_227 (N1722, N763_t1, N1340_t0);
nand NAND2_228 (N1725, N763_t2, N1340_t1);
not NOT1_229 (N1726, N1268_t0);
nand NAND2_230 (N1727, N1493_t0, N1271);
not NOT1_231 (N1728, N1493_t1);
and AND2_232 (N1729, N683_t1, N1268_t1);
nand NAND2_233 (N1730, N1499_t0, N1272);
not NOT1_234 (N1731, N1499_t1);
nand NAND2_235 (N1735, N87_t5, N1264_t1);
not NOT1_236 (N1736, N1273_t0);
not NOT1_237 (N1737, N1276_t0);
nand NAND2_238 (N1738, N1325_t0, N821_t1);
nand NAND2_239 (N1747, N1325_t1, N825_t2);
nand NAND3_240 (N1756, N772_t3, N1279_t0, N798_t2);
nand NAND4_241 (N1761, N772_t4, N786_t3, N798_t3, N1302_t0);
nand NAND2_242 (N1764, N1496_t0, N1339);
not NOT1_243 (N1765, N1496_t1);
nand NAND2_244 (N1766, N1502_t0, N1344);
not NOT1_245 (N1767, N1502_t1);
not NOT1_246 (N1768, N1328_t0);
not NOT1_247 (N1769, N1334_t0);
not NOT1_248 (N1770, N1331_t0);
and AND2_249 (N1787, N845_t0, N1579);
and AND2_250 (N1788, N150_t0, N1580);
and AND2_251 (N1789, N851_t0, N1582);
and AND2_252 (N1790, N159_t0, N1583);
and AND2_253 (N1791, N77_t4, N1584);
and AND2_254 (N1792, N50_t4, N1585);
and AND2_255 (N1793, N858_t0, N1587);
and AND2_256 (N1794, N845_t1, N1588);
and AND2_257 (N1795, N864_t0, N1590);
and AND2_258 (N1796, N851_t1, N1591);
and AND2_259 (N1797, N107_t4, N1593);
and AND2_260 (N1798, N77_t5, N1594);
and AND2_261 (N1799, N116_t3, N1595);
and AND2_262 (N1800, N858_t1, N1596);
and AND2_263 (N1801, N283_t0, N1598);
and AND2_264 (N1802, N864_t1, N1599);
and AND2_265 (N1803, N200_t3, N1363_t0);
and AND2_266 (N1806, N889, N1363_t1);
and AND2_267 (N1809, N890, N1366_t0);
and AND2_268 (N1812, N891, N1366_t1);
nand NAND2_269 (N1815, N1298_t0, N1302_t1);
nand NAND2_270 (N1818, N821_t2, N1302_t2);
nand NAND3_271 (N1821, N772_t5, N1279_t1, N1179);
nand NAND3_272 (N1824, N786_t4, N794_t2, N1298_t1);
nand NAND2_273 (N1833, N786_t5, N1298_t2);
not NOT1_274 (N1842, N1369_t0);
not NOT1_275 (N1843, N1369_t1);
not NOT1_276 (N1844, N1369_t2);
not NOT1_277 (N1845, N1369_t3);
not NOT1_278 (N1846, N1369_t4);
not NOT1_279 (N1847, N1369_t5);
not NOT1_280 (N1848, N1369_t6);
not NOT1_281 (N1849, N1384_t0);
and AND2_282 (N1850, N1384_t1, N896_t8);
not NOT1_283 (N1851, N1384_t2);
and AND2_284 (N1852, N1384_t3, N896_t9);
not NOT1_285 (N1853, N1384_t4);
and AND2_286 (N1854, N1384_t5, N896_t10);
not NOT1_287 (N1855, N1384_t6);
and AND2_288 (N1856, N1384_t7, N896_t11);
not NOT1_289 (N1857, N1384_t8);
and AND2_290 (N1858, N1384_t9, N896_t12);
not NOT1_291 (N1859, N1384_t10);
and AND2_292 (N1860, N1384_t11, N896_t13);
not NOT1_293 (N1861, N1384_t12);
and AND2_294 (N1862, N1384_t13, N896_t14);
not NOT1_295 (N1863, N1384_t14);
and AND2_296 (N1864, N1384_t15, N896_t15);
and AND2_297 (N1869, N1202_t8, N1409_t0);
nor NOR2_298 (N1870, N50_t5, N1409_t1);
not NOT1_299 (N1873, N1306_t0);
and AND2_300 (N1874, N1202_t9, N1409_t2);
nor NOR2_301 (N1875, N58_t6, N1409_t3);
not NOT1_302 (N1878, N1306_t1);
and AND2_303 (N1879, N1202_t10, N1409_t4);
nor NOR2_304 (N1880, N68_t6, N1409_t5);
not NOT1_305 (N1883, N1306_t2);
and AND2_306 (N1884, N1202_t11, N1409_t6);
nor NOR2_307 (N1885, N77_t6, N1409_t7);
not NOT1_308 (N1888, N1306_t3);
and AND2_309 (N1889, N1202_t12, N1409_t8);
nor NOR2_310 (N1890, N87_t6, N1409_t9);
not NOT1_311 (N1893, N1322_t0);
and AND2_312 (N1894, N1202_t13, N1409_t10);
nor NOR2_313 (N1895, N97_t6, N1409_t11);
not NOT1_314 (N1898, N1315_t0);
and AND2_315 (N1899, N1202_t14, N1409_t12);
nor NOR2_316 (N1900, N107_t5, N1409_t13);
not NOT1_317 (N1903, N1315_t1);
and AND2_318 (N1904, N1202_t15, N1409_t14);
nor NOR2_319 (N1905, N116_t4, N1409_t15);
not NOT1_320 (N1908, N1315_t2);
and AND2_321 (N1909, N1452_t0, N213_t1);
nand NAND2_322 (N1912, N1452_t1, N213_t2);
and AND3_323 (N1913, N1452_t2, N213_t3, N343_t1);
nand NAND3_324 (N1917, N1452_t3, N213_t4, N343_t2);
and AND3_325 (N1922, N1452_t4, N213_t5, N343_t3);
nand NAND3_326 (N1926, N1452_t5, N213_t6, N343_t4);
buf BUFF1_327 (N1930, N1464_t0);
nand NAND2_328 (N1933, N1691, N1692);
nand NAND2_329 (N1936, N1693, N1694);
not NOT1_330 (N1939, N1471_t0);
nand NAND2_331 (N1940, N1471_t1, N1474);
not NOT1_332 (N1941, N1475_t0);
not NOT1_333 (N1942, N1478_t0);
not NOT1_334 (N1943, N1481_t0);
not NOT1_335 (N1944, N1484_t0);
not NOT1_336 (N1945, N1487_t0);
not NOT1_337 (N1946, N1490_t0);
not NOT1_338 (N1947, N1714);
nand NAND2_339 (N1960, N953_t1, N1728);
nand NAND2_340 (N1961, N959_t1, N1731);
and AND2_341 (N1966, N1520_t0, N1276_t1);
nand NAND2_342 (N1981, N956_t1, N1765);
nand NAND2_343 (N1982, N962_t1, N1767);
and AND2_344 (N1983, N1067, N1768);
or OR3_345 (N1986, N1581, N1787, N1788);
or OR3_346 (N1987, N1586, N1791, N1792);
or OR3_347 (N1988, N1589, N1793, N1794);
or OR3_348 (N1989, N1592, N1795, N1796);
or OR3_349 (N1990, N1597, N1799, N1800);
or OR3_350 (N1991, N1600, N1801, N1802);
and AND2_351 (N2022, N77_t7, N1849);
and AND2_352 (N2023, N223_t1, N1850);
and AND2_353 (N2024, N87_t7, N1851);
and AND2_354 (N2025, N226_t3, N1852);
and AND2_355 (N2026, N97_t7, N1853);
and AND2_356 (N2027, N232_t3, N1854);
and AND2_357 (N2028, N107_t6, N1855);
and AND2_358 (N2029, N238_t3, N1856);
and AND2_359 (N2030, N116_t5, N1857);
and AND2_360 (N2031, N244_t3, N1858);
and AND2_361 (N2032, N283_t1, N1859);
and AND2_362 (N2033, N250_t4, N1860);
and AND2_363 (N2034, N294_t0, N1861);
and AND2_364 (N2035, N257_t4, N1862);
and AND2_365 (N2036, N303_t0, N1863);
and AND2_366 (N2037, N264_t3, N1864);
buf BUFF1_367 (N2038, N1667_t0);
not NOT1_368 (N2043, N1667_t1);
buf BUFF1_369 (N2052, N1670_t0);
not NOT1_370 (N2057, N1670_t1);
and AND3_371 (N2068, N50_t6, N1197_t0, N1869);
and AND3_372 (N2073, N58_t7, N1197_t1, N1874);
and AND3_373 (N2078, N68_t7, N1197_t2, N1879);
and AND3_374 (N2083, N77_t8, N1197_t3, N1884);
and AND3_375 (N2088, N87_t8, N1219_t0, N1889);
and AND3_376 (N2093, N97_t8, N1219_t1, N1894);
and AND3_377 (N2098, N107_t7, N1219_t2, N1899);
and AND3_378 (N2103, N116_t6, N1219_t3, N1904);
not NOT1_379 (N2121, N1562_t0);
not NOT1_380 (N2122, N1562_t1);
not NOT1_381 (N2123, N1562_t2);
not NOT1_382 (N2124, N1562_t3);
not NOT1_383 (N2125, N1562_t4);
not NOT1_384 (N2126, N1562_t5);
not NOT1_385 (N2127, N1562_t6);
not NOT1_386 (N2128, N1562_t7);
nand NAND2_387 (N2133, N950_t1, N1939);
nand NAND2_388 (N2134, N1478_t1, N1941);
nand NAND2_389 (N2135, N1475_t1, N1942);
nand NAND2_390 (N2136, N1484_t1, N1943);
nand NAND2_391 (N2137, N1481_t1, N1944);
nand NAND2_392 (N2138, N1490_t1, N1945);
nand NAND2_393 (N2139, N1487_t1, N1946);
not NOT1_394 (N2141, N1933_t0);
not NOT1_395 (N2142, N1936_t0);
not NOT1_396 (N2143, N1738_t0);
and AND2_397 (N2144, N1738_t1, N1747_t0);
not NOT1_398 (N2145, N1747_t1);
nand NAND2_399 (N2146, N1727, N1960);
nand NAND2_400 (N2147, N1730, N1961);
and AND4_401 (N2148, N1722_t0, N1267, N665_t1, N58_t8);
not NOT1_402 (N2149, N1738_t2);
and AND2_403 (N2150, N1738_t3, N1747_t2);
not NOT1_404 (N2151, N1747_t3);
not NOT1_405 (N2152, N1738_t4);
not NOT1_406 (N2153, N1747_t4);
and AND2_407 (N2154, N1738_t5, N1747_t5);
not NOT1_408 (N2155, N1738_t6);
not NOT1_409 (N2156, N1747_t6);
and AND2_410 (N2157, N1738_t7, N1747_t7);
buf BUFF1_411 (N2158, N1761_t0);
buf BUFF1_412 (N2175, N1761_t1);
nand NAND2_413 (N2178, N1764, N1981);
nand NAND2_414 (N2179, N1766, N1982);
not NOT1_415 (N2180, N1756_t0);
and AND2_416 (N2181, N1756_t1, N1328_t1);
not NOT1_417 (N2183, N1756_t2);
and AND2_418 (N2184, N1331_t1, N1756_t3);
nand NAND2_419 (N2185, N1358_t0, N1812_t0);
nand NAND2_420 (N2188, N1358_t1, N1809_t0);
nand NAND2_421 (N2191, N1353_t0, N1812_t1);
nand NAND2_422 (N2194, N1353_t1, N1809_t1);
nand NAND2_423 (N2197, N1358_t2, N1806_t0);
nand NAND2_424 (N2200, N1358_t3, N1803_t0);
nand NAND2_425 (N2203, N1353_t2, N1806_t1);
nand NAND2_426 (N2206, N1353_t3, N1803_t1);
not NOT1_427 (N2209, N1815_t0);
not NOT1_428 (N2210, N1818_t0);
and AND2_429 (N2211, N1815_t1, N1818_t1);
buf BUFF1_430 (N2212, N1821_t0);
buf BUFF1_431 (N2221, N1821_t1);
not NOT1_432 (N2230, N1833_t0);
not NOT1_433 (N2231, N1833_t1);
not NOT1_434 (N2232, N1833_t2);
not NOT1_435 (N2233, N1833_t3);
not NOT1_436 (N2234, N1824_t0);
not NOT1_437 (N2235, N1824_t1);
not NOT1_438 (N2236, N1824_t2);
not NOT1_439 (N2237, N1824_t3);
or OR3_440 (N2238, N2022, N1643, N2023);
or OR3_441 (N2239, N2024, N1644, N2025);
or OR3_442 (N2240, N2026, N1645, N2027);
or OR3_443 (N2241, N2028, N1646, N2029);
or OR3_444 (N2242, N2030, N1647, N2031);
or OR3_445 (N2243, N2032, N1648, N2033);
or OR3_446 (N2244, N2034, N1649, N2035);
or OR3_447 (N2245, N2036, N1650, N2037);
and AND2_448 (N2270, N1986, N1673);
and AND2_449 (N2277, N1987, N1675);
and AND2_450 (N2282, N1988, N1676);
and AND2_451 (N2287, N1989, N1677);
and AND2_452 (N2294, N1990, N1679);
and AND2_453 (N2299, N1991, N1680);
buf BUFF1_454 (N2304, N1917_t0);
and AND2_455 (N2307, N1930_t0, N350_t0);
nand NAND2_456 (N2310, N1930_t1, N350_t1);
buf BUFF1_457 (N2313, N1715_t0);
buf BUFF1_458 (N2316, N1718_t0);
buf BUFF1_459 (N2319, N1715_t1);
buf BUFF1_460 (N2322, N1718_t1);
nand NAND2_461 (N2325, N1940, N2133);
nand NAND2_462 (N2328, N2134, N2135);
nand NAND2_463 (N2331, N2136, N2137);
nand NAND2_464 (N2334, N2138, N2139);
nand NAND2_465 (N2341, N1936_t1, N2141);
nand NAND2_466 (N2342, N1933_t1, N2142);
and AND2_467 (N2347, N724_t1, N2144);
and AND3_468 (N2348, N2146, N699_t1, N1726);
and AND2_469 (N2349, N753_t1, N2147);
and AND2_470 (N2350, N2148, N1273_t1);
and AND2_471 (N2351, N736_t2, N2150);
and AND2_472 (N2352, N1735, N2153);
and AND2_473 (N2353, N763_t3, N2154);
and AND2_474 (N2354, N1725, N2156);
and AND2_475 (N2355, N749_t2, N2157);
not NOT1_476 (N2374, N2178);
not NOT1_477 (N2375, N2179);
and AND2_478 (N2376, N1520_t1, N2180);
and AND2_479 (N2379, N1721, N2181);
and AND2_480 (N2398, N665_t2, N2211);
and AND3_481 (N2417, N2057_t0, N226_t4, N1873);
and AND3_482 (N2418, N2057_t1, N274_t0, N1306_t4);
and AND2_483 (N2419, N2052_t0, N2238);
and AND3_484 (N2420, N2057_t2, N232_t4, N1878);
and AND3_485 (N2421, N2057_t3, N274_t1, N1306_t5);
and AND2_486 (N2422, N2052_t1, N2239);
and AND3_487 (N2425, N2057_t4, N238_t4, N1883);
and AND3_488 (N2426, N2057_t5, N274_t2, N1306_t6);
and AND2_489 (N2427, N2052_t2, N2240);
and AND3_490 (N2430, N2057_t6, N244_t4, N1888);
and AND3_491 (N2431, N2057_t7, N274_t3, N1306_t7);
and AND2_492 (N2432, N2052_t3, N2241);
and AND3_493 (N2435, N2043_t0, N250_t5, N1893);
and AND3_494 (N2436, N2043_t1, N274_t4, N1322_t1);
and AND2_495 (N2437, N2038_t0, N2242);
and AND3_496 (N2438, N2043_t2, N257_t5, N1898);
and AND3_497 (N2439, N2043_t3, N274_t5, N1315_t3);
and AND2_498 (N2440, N2038_t1, N2243);
and AND3_499 (N2443, N2043_t4, N264_t4, N1903);
and AND3_500 (N2444, N2043_t5, N274_t6, N1315_t4);
and AND2_501 (N2445, N2038_t2, N2244);
and AND3_502 (N2448, N2043_t6, N270_t2, N1908);
and AND3_503 (N2449, N2043_t7, N274_t7, N1315_t5);
and AND2_504 (N2450, N2038_t3, N2245);
not NOT1_505 (N2467, N2313_t0);
not NOT1_506 (N2468, N2316_t0);
not NOT1_507 (N2469, N2319_t0);
not NOT1_508 (N2470, N2322_t0);
nand NAND2_509 (N2471, N2341, N2342);
not NOT1_510 (N2474, N2325_t0);
not NOT1_511 (N2475, N2328_t0);
not NOT1_512 (N2476, N2331_t0);
not NOT1_513 (N2477, N2334_t0);
or OR2_514 (N2478, N2348, N1729);
not NOT1_515 (N2481, N2175_t0);
and AND2_516 (N2482, N2175_t1, N1334_t1);
and AND2_517 (N2483, N2349, N2183);
and AND2_518 (N2486, N2374, N1346);
and AND2_519 (N2487, N2375, N1350);
buf BUFF1_520 (N2488, N2185_t0);
buf BUFF1_521 (N2497, N2188_t0);
buf BUFF1_522 (N2506, N2191_t0);
buf BUFF1_523 (N2515, N2194_t0);
buf BUFF1_524 (N2524, N2197_t0);
buf BUFF1_525 (N2533, N2200_t0);
buf BUFF1_526 (N2542, N2203_t0);
buf BUFF1_527 (N2551, N2206_t0);
buf BUFF1_528 (N2560, N2185_t1);
buf BUFF1_529 (N2569, N2188_t1);
buf BUFF1_530 (N2578, N2191_t1);
buf BUFF1_531 (N2587, N2194_t1);
buf BUFF1_532 (N2596, N2197_t1);
buf BUFF1_533 (N2605, N2200_t1);
buf BUFF1_534 (N2614, N2203_t1);
buf BUFF1_535 (N2623, N2206_t1);
not NOT1_536 (N2632, N2212_t0);
and AND2_537 (N2633, N2212_t1, N1833_t4);
not NOT1_538 (N2634, N2212_t2);
and AND2_539 (N2635, N2212_t3, N1833_t5);
not NOT1_540 (N2636, N2212_t4);
and AND2_541 (N2637, N2212_t5, N1833_t6);
not NOT1_542 (N2638, N2212_t6);
and AND2_543 (N2639, N2212_t7, N1833_t7);
not NOT1_544 (N2640, N2221_t0);
and AND2_545 (N2641, N2221_t1, N1824_t4);
not NOT1_546 (N2642, N2221_t2);
and AND2_547 (N2643, N2221_t3, N1824_t5);
not NOT1_548 (N2644, N2221_t4);
and AND2_549 (N2645, N2221_t5, N1824_t6);
not NOT1_550 (N2646, N2221_t6);
and AND2_551 (N2647, N2221_t7, N1824_t7);
or OR3_552 (N2648, N2270_t0, N1870_t0, N2068_t0);
nor NOR3_553 (N2652, N2270_t1, N1870_t1, N2068_t1);
or OR3_554 (N2656, N2417, N2418, N2419);
or OR3_555 (N2659, N2420, N2421, N2422);
or OR3_556 (N2662, N2277_t0, N1880_t0, N2078_t0);
nor NOR3_557 (N2666, N2277_t1, N1880_t1, N2078_t1);
or OR3_558 (N2670, N2425, N2426, N2427);
or OR3_559 (N2673, N2282_t0, N1885_t0, N2083_t0);
nor NOR3_560 (N2677, N2282_t1, N1885_t1, N2083_t1);
or OR3_561 (N2681, N2430, N2431, N2432);
or OR3_562 (N2684, N2287_t0, N1890_t0, N2088_t0);
nor NOR3_563 (N2688, N2287_t1, N1890_t1, N2088_t1);
or OR3_564 (N2692, N2435, N2436, N2437);
or OR3_565 (N2697, N2438, N2439, N2440);
or OR3_566 (N2702, N2294_t0, N1900_t0, N2098_t0);
nor NOR3_567 (N2706, N2294_t1, N1900_t1, N2098_t1);
or OR3_568 (N2710, N2443, N2444, N2445);
or OR3_569 (N2715, N2299_t0, N1905_t0, N2103_t0);
nor NOR3_570 (N2719, N2299_t1, N1905_t1, N2103_t1);
or OR3_571 (N2723, N2448, N2449, N2450);
not NOT1_572 (N2728, N2304_t0);
not NOT1_573 (N2729, N2158_t0);
and AND2_574 (N2730, N1562_t8, N2158_t1);
not NOT1_575 (N2731, N2158_t2);
and AND2_576 (N2732, N1562_t9, N2158_t3);
not NOT1_577 (N2733, N2158_t4);
and AND2_578 (N2734, N1562_t10, N2158_t5);
not NOT1_579 (N2735, N2158_t6);
and AND2_580 (N2736, N1562_t11, N2158_t7);
not NOT1_581 (N2737, N2158_t8);
and AND2_582 (N2738, N1562_t12, N2158_t9);
not NOT1_583 (N2739, N2158_t10);
and AND2_584 (N2740, N1562_t13, N2158_t11);
not NOT1_585 (N2741, N2158_t12);
and AND2_586 (N2742, N1562_t14, N2158_t13);
not NOT1_587 (N2743, N2158_t14);
and AND2_588 (N2744, N1562_t15, N2158_t15);
or OR3_589 (N2745, N2376_t0, N1983_t0, N2379_t0);
nor NOR3_590 (N2746, N2376_t1, N1983_t1, N2379_t1);
nand NAND2_591 (N2748, N2316_t1, N2467);
nand NAND2_592 (N2749, N2313_t1, N2468);
nand NAND2_593 (N2750, N2322_t1, N2469);
nand NAND2_594 (N2751, N2319_t1, N2470);
nand NAND2_595 (N2754, N2328_t1, N2474);
nand NAND2_596 (N2755, N2325_t1, N2475);
nand NAND2_597 (N2756, N2334_t1, N2476);
nand NAND2_598 (N2757, N2331_t1, N2477);
and AND2_599 (N2758, N1520_t2, N2481);
and AND2_600 (N2761, N1722_t1, N2482);
and AND2_601 (N2764, N2478, N1770);
or OR3_602 (N2768, N2486, N1789, N1790);
or OR3_603 (N2769, N2487, N1797, N1798);
and AND2_604 (N2898, N665_t3, N2633);
and AND2_605 (N2899, N679_t2, N2635);
and AND2_606 (N2900, N686_t2, N2637);
and AND2_607 (N2901, N702_t2, N2639);
not NOT1_608 (N2962, N2746);
nand NAND2_609 (N2966, N2748, N2749);
nand NAND2_610 (N2967, N2750, N2751);
buf BUFF1_611 (N2970, N2471_t0);
nand NAND2_612 (N2973, N2754, N2755);
nand NAND2_613 (N2977, N2756, N2757);
and AND2_614 (N2980, N2471_t1, N2143);
not NOT1_615 (N2984, N2488_t0);
not NOT1_616 (N2985, N2497_t0);
not NOT1_617 (N2986, N2506_t0);
not NOT1_618 (N2987, N2515_t0);
not NOT1_619 (N2988, N2524_t0);
not NOT1_620 (N2989, N2533_t0);
not NOT1_621 (N2990, N2542_t0);
not NOT1_622 (N2991, N2551_t0);
not NOT1_623 (N2992, N2488_t1);
not NOT1_624 (N2993, N2497_t1);
not NOT1_625 (N2994, N2506_t1);
not NOT1_626 (N2995, N2515_t1);
not NOT1_627 (N2996, N2524_t1);
not NOT1_628 (N2997, N2533_t1);
not NOT1_629 (N2998, N2542_t1);
not NOT1_630 (N2999, N2551_t1);
not NOT1_631 (N3000, N2488_t2);
not NOT1_632 (N3001, N2497_t2);
not NOT1_633 (N3002, N2506_t2);
not NOT1_634 (N3003, N2515_t2);
not NOT1_635 (N3004, N2524_t2);
not NOT1_636 (N3005, N2533_t2);
not NOT1_637 (N3006, N2542_t2);
not NOT1_638 (N3007, N2551_t2);
not NOT1_639 (N3008, N2488_t3);
not NOT1_640 (N3009, N2497_t3);
not NOT1_641 (N3010, N2506_t3);
not NOT1_642 (N3011, N2515_t3);
not NOT1_643 (N3012, N2524_t3);
not NOT1_644 (N3013, N2533_t3);
not NOT1_645 (N3014, N2542_t3);
not NOT1_646 (N3015, N2551_t3);
not NOT1_647 (N3016, N2488_t4);
not NOT1_648 (N3017, N2497_t4);
not NOT1_649 (N3018, N2506_t4);
not NOT1_650 (N3019, N2515_t4);
not NOT1_651 (N3020, N2524_t4);
not NOT1_652 (N3021, N2533_t4);
not NOT1_653 (N3022, N2542_t4);
not NOT1_654 (N3023, N2551_t4);
not NOT1_655 (N3024, N2488_t5);
not NOT1_656 (N3025, N2497_t5);
not NOT1_657 (N3026, N2506_t5);
not NOT1_658 (N3027, N2515_t5);
not NOT1_659 (N3028, N2524_t5);
not NOT1_660 (N3029, N2533_t5);
not NOT1_661 (N3030, N2542_t5);
not NOT1_662 (N3031, N2551_t5);
not NOT1_663 (N3032, N2488_t6);
not NOT1_664 (N3033, N2497_t6);
not NOT1_665 (N3034, N2506_t6);
not NOT1_666 (N3035, N2515_t6);
not NOT1_667 (N3036, N2524_t6);
not NOT1_668 (N3037, N2533_t6);
not NOT1_669 (N3038, N2542_t6);
not NOT1_670 (N3039, N2551_t6);
not NOT1_671 (N3040, N2488_t7);
not NOT1_672 (N3041, N2497_t7);
not NOT1_673 (N3042, N2506_t7);
not NOT1_674 (N3043, N2515_t7);
not NOT1_675 (N3044, N2524_t7);
not NOT1_676 (N3045, N2533_t7);
not NOT1_677 (N3046, N2542_t7);
not NOT1_678 (N3047, N2551_t7);
not NOT1_679 (N3048, N2560_t0);
not NOT1_680 (N3049, N2569_t0);
not NOT1_681 (N3050, N2578_t0);
not NOT1_682 (N3051, N2587_t0);
not NOT1_683 (N3052, N2596_t0);
not NOT1_684 (N3053, N2605_t0);
not NOT1_685 (N3054, N2614_t0);
not NOT1_686 (N3055, N2623_t0);
not NOT1_687 (N3056, N2560_t1);
not NOT1_688 (N3057, N2569_t1);
not NOT1_689 (N3058, N2578_t1);
not NOT1_690 (N3059, N2587_t1);
not NOT1_691 (N3060, N2596_t1);
not NOT1_692 (N3061, N2605_t1);
not NOT1_693 (N3062, N2614_t1);
not NOT1_694 (N3063, N2623_t1);
not NOT1_695 (N3064, N2560_t2);
not NOT1_696 (N3065, N2569_t2);
not NOT1_697 (N3066, N2578_t2);
not NOT1_698 (N3067, N2587_t2);
not NOT1_699 (N3068, N2596_t2);
not NOT1_700 (N3069, N2605_t2);
not NOT1_701 (N3070, N2614_t2);
not NOT1_702 (N3071, N2623_t2);
not NOT1_703 (N3072, N2560_t3);
not NOT1_704 (N3073, N2569_t3);
not NOT1_705 (N3074, N2578_t3);
not NOT1_706 (N3075, N2587_t3);
not NOT1_707 (N3076, N2596_t3);
not NOT1_708 (N3077, N2605_t3);
not NOT1_709 (N3078, N2614_t3);
not NOT1_710 (N3079, N2623_t3);
not NOT1_711 (N3080, N2560_t4);
not NOT1_712 (N3081, N2569_t4);
not NOT1_713 (N3082, N2578_t4);
not NOT1_714 (N3083, N2587_t4);
not NOT1_715 (N3084, N2596_t4);
not NOT1_716 (N3085, N2605_t4);
not NOT1_717 (N3086, N2614_t4);
not NOT1_718 (N3087, N2623_t4);
not NOT1_719 (N3088, N2560_t5);
not NOT1_720 (N3089, N2569_t5);
not NOT1_721 (N3090, N2578_t5);
not NOT1_722 (N3091, N2587_t5);
not NOT1_723 (N3092, N2596_t5);
not NOT1_724 (N3093, N2605_t5);
not NOT1_725 (N3094, N2614_t5);
not NOT1_726 (N3095, N2623_t5);
not NOT1_727 (N3096, N2560_t6);
not NOT1_728 (N3097, N2569_t6);
not NOT1_729 (N3098, N2578_t6);
not NOT1_730 (N3099, N2587_t6);
not NOT1_731 (N3100, N2596_t6);
not NOT1_732 (N3101, N2605_t6);
not NOT1_733 (N3102, N2614_t6);
not NOT1_734 (N3103, N2623_t6);
not NOT1_735 (N3104, N2560_t7);
not NOT1_736 (N3105, N2569_t7);
not NOT1_737 (N3106, N2578_t7);
not NOT1_738 (N3107, N2587_t7);
not NOT1_739 (N3108, N2596_t7);
not NOT1_740 (N3109, N2605_t7);
not NOT1_741 (N3110, N2614_t7);
not NOT1_742 (N3111, N2623_t7);
buf BUFF1_743 (N3112, N2656_t0);
not NOT1_744 (N3115, N2656_t1);
not NOT1_745 (N3118, N2652_t0);
and AND2_746 (N3119, N2768, N1674);
buf BUFF1_747 (N3122, N2659_t0);
not NOT1_748 (N3125, N2659_t1);
buf BUFF1_749 (N3128, N2670_t0);
not NOT1_750 (N3131, N2670_t1);
not NOT1_751 (N3134, N2666_t0);
buf BUFF1_752 (N3135, N2681_t0);
not NOT1_753 (N3138, N2681_t1);
not NOT1_754 (N3141, N2677_t0);
buf BUFF1_755 (N3142, N2692_t0);
not NOT1_756 (N3145, N2692_t1);
not NOT1_757 (N3148, N2688_t0);
and AND2_758 (N3149, N2769, N1678);
buf BUFF1_759 (N3152, N2697_t0);
not NOT1_760 (N3155, N2697_t1);
buf BUFF1_761 (N3158, N2710_t0);
not NOT1_762 (N3161, N2710_t1);
not NOT1_763 (N3164, N2706_t0);
buf BUFF1_764 (N3165, N2723_t0);
not NOT1_765 (N3168, N2723_t1);
not NOT1_766 (N3171, N2719_t0);
and AND2_767 (N3172, N1909_t0, N2648_t0);
and AND2_768 (N3175, N1913_t0, N2662_t0);
and AND2_769 (N3178, N1913_t1, N2673_t0);
and AND2_770 (N3181, N1913_t2, N2684_t0);
and AND2_771 (N3184, N1922_t0, N2702_t0);
and AND2_772 (N3187, N1922_t1, N2715_t0);
not NOT1_773 (N3190, N2692_t2);
not NOT1_774 (N3191, N2697_t2);
not NOT1_775 (N3192, N2710_t2);
not NOT1_776 (N3193, N2723_t2);
and AND5_777 (N3194, N2692_t3, N2697_t3, N2710_t3, N2723_t3, N1459);
nand NAND2_778 (N3195, N2745, N2962);
not NOT1_779 (N3196, N2966);
or OR3_780 (N3206, N2980, N2145, N2347);
and AND2_781 (N3207, N124_t, N2984);
and AND2_782 (N3208, N159_t1, N2985);
and AND2_783 (N3209, N150_t1, N2986);
and AND2_784 (N3210, N143_t0, N2987);
and AND2_785 (N3211, N137_t0, N2988);
and AND2_786 (N3212, N132_t0, N2989);
and AND2_787 (N3213, N128_t0, N2990);
and AND2_788 (N3214, N125_t0, N2991);
and AND2_789 (N3215, N125_t1, N2992);
and AND2_790 (N3216, N655_t2, N2993);
and AND2_791 (N3217, N159_t2, N2994);
and AND2_792 (N3218, N150_t2, N2995);
and AND2_793 (N3219, N143_t1, N2996);
and AND2_794 (N3220, N137_t1, N2997);
and AND2_795 (N3221, N132_t1, N2998);
and AND2_796 (N3222, N128_t1, N2999);
and AND2_797 (N3223, N128_t2, N3000);
and AND2_798 (N3224, N670_t1, N3001);
and AND2_799 (N3225, N655_t3, N3002);
and AND2_800 (N3226, N159_t3, N3003);
and AND2_801 (N3227, N150_t3, N3004);
and AND2_802 (N3228, N143_t2, N3005);
and AND2_803 (N3229, N137_t2, N3006);
and AND2_804 (N3230, N132_t2, N3007);
and AND2_805 (N3231, N132_t3, N3008);
and AND2_806 (N3232, N690_t1, N3009);
and AND2_807 (N3233, N670_t2, N3010);
and AND2_808 (N3234, N655_t4, N3011);
and AND2_809 (N3235, N159_t4, N3012);
and AND2_810 (N3236, N150_t4, N3013);
and AND2_811 (N3237, N143_t3, N3014);
and AND2_812 (N3238, N137_t3, N3015);
and AND2_813 (N3239, N137_t4, N3016);
and AND2_814 (N3240, N706_t1, N3017);
and AND2_815 (N3241, N690_t2, N3018);
and AND2_816 (N3242, N670_t3, N3019);
and AND2_817 (N3243, N655_t5, N3020);
and AND2_818 (N3244, N159_t5, N3021);
and AND2_819 (N3245, N150_t5, N3022);
and AND2_820 (N3246, N143_t4, N3023);
and AND2_821 (N3247, N143_t5, N3024);
and AND2_822 (N3248, N715_t1, N3025);
and AND2_823 (N3249, N706_t2, N3026);
and AND2_824 (N3250, N690_t3, N3027);
and AND2_825 (N3251, N670_t4, N3028);
and AND2_826 (N3252, N655_t6, N3029);
and AND2_827 (N3253, N159_t6, N3030);
and AND2_828 (N3254, N150_t6, N3031);
and AND2_829 (N3255, N150_t7, N3032);
and AND2_830 (N3256, N727_t1, N3033);
and AND2_831 (N3257, N715_t2, N3034);
and AND2_832 (N3258, N706_t3, N3035);
and AND2_833 (N3259, N690_t4, N3036);
and AND2_834 (N3260, N670_t5, N3037);
and AND2_835 (N3261, N655_t7, N3038);
and AND2_836 (N3262, N159_t7, N3039);
and AND2_837 (N3263, N159_t8, N3040);
and AND2_838 (N3264, N740_t1, N3041);
and AND2_839 (N3265, N727_t2, N3042);
and AND2_840 (N3266, N715_t3, N3043);
and AND2_841 (N3267, N706_t4, N3044);
and AND2_842 (N3268, N690_t5, N3045);
and AND2_843 (N3269, N670_t6, N3046);
and AND2_844 (N3270, N655_t8, N3047);
and AND2_845 (N3271, N283_t2, N3048);
and AND2_846 (N3272, N670_t7, N3049);
and AND2_847 (N3273, N690_t6, N3050);
and AND2_848 (N3274, N706_t5, N3051);
and AND2_849 (N3275, N715_t4, N3052);
and AND2_850 (N3276, N727_t3, N3053);
and AND2_851 (N3277, N740_t2, N3054);
and AND2_852 (N3278, N753_t2, N3055);
and AND2_853 (N3279, N294_t1, N3056);
and AND2_854 (N3280, N690_t7, N3057);
and AND2_855 (N3281, N706_t6, N3058);
and AND2_856 (N3282, N715_t5, N3059);
and AND2_857 (N3283, N727_t4, N3060);
and AND2_858 (N3284, N740_t3, N3061);
and AND2_859 (N3285, N753_t3, N3062);
and AND2_860 (N3286, N283_t3, N3063);
and AND2_861 (N3287, N303_t1, N3064);
and AND2_862 (N3288, N706_t7, N3065);
and AND2_863 (N3289, N715_t6, N3066);
and AND2_864 (N3290, N727_t5, N3067);
and AND2_865 (N3291, N740_t4, N3068);
and AND2_866 (N3292, N753_t4, N3069);
and AND2_867 (N3293, N283_t4, N3070);
and AND2_868 (N3294, N294_t2, N3071);
and AND2_869 (N3295, N311_t0, N3072);
and AND2_870 (N3296, N715_t7, N3073);
and AND2_871 (N3297, N727_t6, N3074);
and AND2_872 (N3298, N740_t5, N3075);
and AND2_873 (N3299, N753_t5, N3076);
and AND2_874 (N3300, N283_t5, N3077);
and AND2_875 (N3301, N294_t3, N3078);
and AND2_876 (N3302, N303_t2, N3079);
and AND2_877 (N3303, N317_t0, N3080);
and AND2_878 (N3304, N727_t7, N3081);
and AND2_879 (N3305, N740_t6, N3082);
and AND2_880 (N3306, N753_t6, N3083);
and AND2_881 (N3307, N283_t6, N3084);
and AND2_882 (N3308, N294_t4, N3085);
and AND2_883 (N3309, N303_t3, N3086);
and AND2_884 (N3310, N311_t1, N3087);
and AND2_885 (N3311, N322_t0, N3088);
and AND2_886 (N3312, N740_t7, N3089);
and AND2_887 (N3313, N753_t7, N3090);
and AND2_888 (N3314, N283_t7, N3091);
and AND2_889 (N3315, N294_t5, N3092);
and AND2_890 (N3316, N303_t4, N3093);
and AND2_891 (N3317, N311_t2, N3094);
and AND2_892 (N3318, N317_t1, N3095);
and AND2_893 (N3319, N326_t0, N3096);
and AND2_894 (N3320, N753_t8, N3097);
and AND2_895 (N3321, N283_t8, N3098);
and AND2_896 (N3322, N294_t6, N3099);
and AND2_897 (N3323, N303_t5, N3100);
and AND2_898 (N3324, N311_t3, N3101);
and AND2_899 (N3325, N317_t2, N3102);
and AND2_900 (N3326, N322_t1, N3103);
and AND2_901 (N3327, N329_t, N3104);
and AND2_902 (N3328, N283_t9, N3105);
and AND2_903 (N3329, N294_t7, N3106);
and AND2_904 (N3330, N303_t6, N3107);
and AND2_905 (N3331, N311_t4, N3108);
and AND2_906 (N3332, N317_t3, N3109);
and AND2_907 (N3333, N322_t2, N3110);
and AND2_908 (N3334, N326_t1, N3111);
and AND5_909 (N3383, N3190, N3191, N3192, N3193, N917_t1);
buf BUFF1_910 (N3384, N2977_t0);
and AND2_911 (N3387, N3196, N1736);
and AND2_912 (N3388, N2977_t1, N2149);
and AND2_913 (N3389, N2973_t0, N1737);
nor NOR8_914 (N3390, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214);
nor NOR8_915 (N3391, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222);
nor NOR8_916 (N3392, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230);
nor NOR8_917 (N3393, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238);
nor NOR8_918 (N3394, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246);
nor NOR8_919 (N3395, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254);
nor NOR8_920 (N3396, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262);
nor NOR8_921 (N3397, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270);
nor NOR8_922 (N3398, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278);
nor NOR8_923 (N3399, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286);
nor NOR8_924 (N3400, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294);
nor NOR8_925 (N3401, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302);
nor NOR8_926 (N3402, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310);
nor NOR8_927 (N3403, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318);
nor NOR8_928 (N3404, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326);
nor NOR8_929 (N3405, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334);
and AND2_930 (N3406, N3206, N2641);
and AND3_931 (N3407, N169_t1, N2648_t1, N3112_t0);
and AND3_932 (N3410, N179_t2, N2648_t2, N3115_t0);
and AND3_933 (N3413, N190_t1, N2652_t1, N3115_t1);
and AND3_934 (N3414, N200_t4, N2652_t2, N3112_t1);
or OR3_935 (N3415, N3119_t0, N1875_t0, N2073_t0);
nor NOR3_936 (N3419, N3119_t1, N1875_t1, N2073_t1);
and AND3_937 (N3423, N169_t2, N2662_t1, N3128_t0);
and AND3_938 (N3426, N179_t3, N2662_t2, N3131_t0);
and AND3_939 (N3429, N190_t2, N2666_t1, N3131_t1);
and AND3_940 (N3430, N200_t5, N2666_t2, N3128_t1);
and AND3_941 (N3431, N169_t3, N2673_t1, N3135_t0);
and AND3_942 (N3434, N179_t4, N2673_t2, N3138_t0);
and AND3_943 (N3437, N190_t3, N2677_t1, N3138_t1);
and AND3_944 (N3438, N200_t6, N2677_t2, N3135_t1);
and AND3_945 (N3439, N169_t4, N2684_t1, N3142_t0);
and AND3_946 (N3442, N179_t5, N2684_t2, N3145_t0);
and AND3_947 (N3445, N190_t4, N2688_t1, N3145_t1);
and AND3_948 (N3446, N200_t7, N2688_t2, N3142_t1);
or OR3_949 (N3447, N3149_t0, N1895_t0, N2093_t0);
nor NOR3_950 (N3451, N3149_t1, N1895_t1, N2093_t1);
and AND3_951 (N3455, N169_t5, N2702_t1, N3158_t0);
and AND3_952 (N3458, N179_t6, N2702_t2, N3161_t0);
and AND3_953 (N3461, N190_t5, N2706_t1, N3161_t1);
and AND3_954 (N3462, N200_t8, N2706_t2, N3158_t1);
and AND3_955 (N3463, N169_t6, N2715_t1, N3165_t0);
and AND3_956 (N3466, N179_t7, N2715_t2, N3168_t0);
and AND3_957 (N3469, N190_t6, N2719_t1, N3168_t1);
and AND3_958 (N3470, N200_t9, N2719_t2, N3165_t1);
or OR2_959 (N3471, N3194, N3383);
buf BUFF1_960 (N3472, N2967_t0);
buf BUFF1_961 (N3475, N2970_t0);
buf BUFF1_962 (N3478, N2967_t1);
buf BUFF1_963 (N3481, N2970_t1);
buf BUFF1_964 (N3484, N2973_t1);
buf BUFF1_965 (N3487, N2973_t2);
buf BUFF1_966 (N3490, N3172_t0);
buf BUFF1_967 (N3493, N3172_t1);
buf BUFF1_968 (N3496, N3175_t0);
buf BUFF1_969 (N3499, N3175_t1);
buf BUFF1_970 (N3502, N3178_t0);
buf BUFF1_971 (N3505, N3178_t1);
buf BUFF1_972 (N3508, N3181_t0);
buf BUFF1_973 (N3511, N3181_t1);
buf BUFF1_974 (N3514, N3184_t0);
buf BUFF1_975 (N3517, N3184_t1);
buf BUFF1_976 (N3520, N3187_t0);
buf BUFF1_977 (N3523, N3187_t1);
nor NOR2_978 (N3534, N3387, N2350);
or OR3_979 (N3535, N3388, N2151, N2351);
nor NOR2_980 (N3536, N3389, N1966);
and AND2_981 (N3537, N3390, N2209);
and AND2_982 (N3538, N3398, N2210);
and AND2_983 (N3539, N3391, N1842);
and AND2_984 (N3540, N3399, N1369_t7);
and AND2_985 (N3541, N3392, N1843);
and AND2_986 (N3542, N3400, N1369_t8);
and AND2_987 (N3543, N3393, N1844);
and AND2_988 (N3544, N3401, N1369_t9);
and AND2_989 (N3545, N3394, N1845);
and AND2_990 (N3546, N3402, N1369_t10);
and AND2_991 (N3547, N3395, N1846);
and AND2_992 (N3548, N3403, N1369_t11);
and AND2_993 (N3549, N3396, N1847);
and AND2_994 (N3550, N3404, N1369_t12);
and AND2_995 (N3551, N3397, N1848);
and AND2_996 (N3552, N3405, N1369_t13);
or OR3_997 (N3557, N3413, N3414, N3118);
or OR3_998 (N3568, N3429, N3430, N3134);
or OR3_999 (N3573, N3437, N3438, N3141);
or OR3_1000 (N3578, N3445, N3446, N3148);
or OR3_1001 (N3589, N3461, N3462, N3164);
or OR3_1002 (N3594, N3469, N3470, N3171);
and AND2_1003 (N3605, N3471, N2728);
not NOT1_1004 (N3626, N3478_t0);
not NOT1_1005 (N3627, N3481_t0);
not NOT1_1006 (N3628, N3487_t0);
not NOT1_1007 (N3629, N3484_t0);
not NOT1_1008 (N3630, N3472_t0);
not NOT1_1009 (N3631, N3475_t0);
and AND2_1010 (N3632, N3536, N2152);
and AND2_1011 (N3633, N3534, N2155);
or OR3_1012 (N3634, N3537, N3538, N2398);
or OR2_1013 (N3635, N3539, N3540);
or OR2_1014 (N3636, N3541, N3542);
or OR2_1015 (N3637, N3543, N3544);
or OR2_1016 (N3638, N3545, N3546);
or OR2_1017 (N3639, N3547, N3548);
or OR2_1018 (N3640, N3549, N3550);
or OR2_1019 (N3641, N3551, N3552);
and AND2_1020 (N3642, N3535, N2643);
or OR2_1021 (N3643, N3407_t0, N3410_t0);
nor NOR2_1022 (N3644, N3407_t1, N3410_t1);
and AND3_1023 (N3645, N169_t7, N3415_t0, N3122_t0);
and AND3_1024 (N3648, N179_t8, N3415_t1, N3125_t0);
and AND3_1025 (N3651, N190_t7, N3419_t0, N3125_t1);
and AND3_1026 (N3652, N200_t10, N3419_t1, N3122_t1);
not NOT1_1027 (N3653, N3419_t2);
or OR2_1028 (N3654, N3423_t0, N3426_t0);
nor NOR2_1029 (N3657, N3423_t1, N3426_t1);
or OR2_1030 (N3658, N3431_t0, N3434_t0);
nor NOR2_1031 (N3661, N3431_t1, N3434_t1);
or OR2_1032 (N3662, N3439_t0, N3442_t0);
nor NOR2_1033 (N3663, N3439_t1, N3442_t1);
and AND3_1034 (N3664, N169_t8, N3447_t0, N3152_t0);
and AND3_1035 (N3667, N179_t9, N3447_t1, N3155_t0);
and AND3_1036 (N3670, N190_t8, N3451_t0, N3155_t1);
and AND3_1037 (N3671, N200_t11, N3451_t1, N3152_t1);
not NOT1_1038 (N3672, N3451_t2);
or OR2_1039 (N3673, N3455_t0, N3458_t0);
nor NOR2_1040 (N3676, N3455_t1, N3458_t1);
or OR2_1041 (N3677, N3463_t0, N3466_t0);
nor NOR2_1042 (N3680, N3463_t1, N3466_t1);
not NOT1_1043 (N3681, N3493_t0);
and AND2_1044 (N3682, N1909_t1, N3415_t2);
not NOT1_1045 (N3685, N3496_t0);
not NOT1_1046 (N3686, N3499_t0);
not NOT1_1047 (N3687, N3502_t0);
not NOT1_1048 (N3688, N3505_t0);
not NOT1_1049 (N3689, N3511_t0);
and AND2_1050 (N3690, N1922_t2, N3447_t2);
not NOT1_1051 (N3693, N3517_t0);
not NOT1_1052 (N3694, N3520_t0);
not NOT1_1053 (N3695, N3523_t0);
not NOT1_1054 (N3696, N3514_t0);
buf BUFF1_1055 (N3697, N3384_t0);
buf BUFF1_1056 (N3700, N3384_t1);
not NOT1_1057 (N3703, N3490_t0);
not NOT1_1058 (N3704, N3508_t0);
nand NAND2_1059 (N3705, N3475_t1, N3630);
nand NAND2_1060 (N3706, N3472_t1, N3631);
nand NAND2_1061 (N3707, N3481_t1, N3626);
nand NAND2_1062 (N3708, N3478_t1, N3627);
or OR3_1063 (N3711, N3632, N2352, N2353);
or OR3_1064 (N3712, N3633, N2354, N2355);
and AND2_1065 (N3713, N3634, N2632);
and AND2_1066 (N3714, N3635, N2634);
and AND2_1067 (N3715, N3636, N2636);
and AND2_1068 (N3716, N3637, N2638);
and AND2_1069 (N3717, N3638, N2640);
and AND2_1070 (N3718, N3639, N2642);
and AND2_1071 (N3719, N3640, N2644);
and AND2_1072 (N3720, N3641, N2646);
and AND2_1073 (N3721, N3644, N3557);
or OR3_1074 (N3731, N3651, N3652, N3653);
and AND2_1075 (N3734, N3657, N3568);
and AND2_1076 (N3740, N3661, N3573);
and AND2_1077 (N3743, N3663, N3578);
or OR3_1078 (N3753, N3670, N3671, N3672);
and AND2_1079 (N3756, N3676, N3589);
and AND2_1080 (N3762, N3680, N3594);
not NOT1_1081 (N3765, N3643);
not NOT1_1082 (N3766, N3662);
nand NAND2_1083 (N3773, N3705, N3706);
nand NAND2_1084 (N3774, N3707, N3708);
nand NAND2_1085 (N3775, N3700_t0, N3628);
not NOT1_1086 (N3776, N3700_t1);
nand NAND2_1087 (N3777, N3697_t0, N3629);
not NOT1_1088 (N3778, N3697_t1);
and AND2_1089 (N3779, N3712, N2645);
and AND2_1090 (N3780, N3711, N2647);
or OR2_1091 (N3786, N3645_t0, N3648_t0);
nor NOR2_1092 (N3789, N3645_t1, N3648_t1);
or OR2_1093 (N3800, N3664_t0, N3667_t0);
nor NOR2_1094 (N3803, N3664_t1, N3667_t1);
and AND2_1095 (N3809, N3654_t0, N1917_t1);
and AND2_1096 (N3812, N3658_t0, N1917_t2);
and AND2_1097 (N3815, N3673_t0, N1926_t0);
and AND2_1098 (N3818, N3677_t0, N1926_t1);
buf BUFF1_1099 (N3821, N3682_t0);
buf BUFF1_1100 (N3824, N3682_t1);
buf BUFF1_1101 (N3827, N3690_t0);
buf BUFF1_1102 (N3830, N3690_t1);
nand NAND2_1103 (N3833, N3773, N3774);
nand NAND2_1104 (N3834, N3487_t1, N3776);
nand NAND2_1105 (N3835, N3484_t1, N3778);
and AND2_1106 (N3838, N3789, N3731);
and AND2_1107 (N3845, N3803, N3753);
buf BUFF1_1108 (N3850, N3721_t0);
buf BUFF1_1109 (N3855, N3734_t0);
buf BUFF1_1110 (N3858, N3740_t0);
buf BUFF1_1111 (N3861, N3743_t0);
buf BUFF1_1112 (N3865, N3756_t0);
buf BUFF1_1113 (N3868, N3762_t0);
nand NAND2_1114 (N3884, N3775, N3834);
nand NAND2_1115 (N3885, N3777, N3835);
nand NAND2_1116 (N3894, N3721_t1, N3786_t0);
nand NAND2_1117 (N3895, N3743_t1, N3800_t0);
not NOT1_1118 (N3898, N3821_t0);
not NOT1_1119 (N3899, N3824_t0);
not NOT1_1120 (N3906, N3830_t0);
not NOT1_1121 (N3911, N3827_t0);
and AND2_1122 (N3912, N3786_t1, N1912);
buf BUFF1_1123 (N3913, N3812_t0);
and AND2_1124 (N3916, N3800_t1, N1917_t3);
buf BUFF1_1125 (N3917, N3818_t0);
not NOT1_1126 (N3920, N3809_t0);
buf BUFF1_1127 (N3921, N3818_t1);
not NOT1_1128 (N3924, N3884);
not NOT1_1129 (N3925, N3885);
and AND4_1130 (N3926, N3721_t2, N3838_t0, N3734_t1, N3740_t1);
nand NAND3_1131 (N3930, N3721_t3, N3838_t1, N3654_t1);
nand NAND4_1132 (N3931, N3658_t1, N3838_t2, N3734_t2, N3721_t4);
and AND4_1133 (N3932, N3743_t2, N3845_t0, N3756_t1, N3762_t1);
nand NAND3_1134 (N3935, N3743_t3, N3845_t1, N3673_t1);
nand NAND4_1135 (N3936, N3677_t1, N3845_t2, N3756_t2, N3743_t4);
buf BUFF1_1136 (N3937, N3838_t3);
buf BUFF1_1137 (N3940, N3845_t3);
not NOT1_1138 (N3947, N3912);
not NOT1_1139 (N3948, N3916);
buf BUFF1_1140 (N3950, N3850_t0);
buf BUFF1_1141 (N3953, N3850_t1);
buf BUFF1_1142 (N3956, N3855_t0);
buf BUFF1_1143 (N3959, N3855_t1);
buf BUFF1_1144 (N3962, N3858_t0);
buf BUFF1_1145 (N3965, N3858_t1);
buf BUFF1_1146 (N3968, N3861_t0);
buf BUFF1_1147 (N3971, N3861_t1);
buf BUFF1_1148 (N3974, N3865_t0);
buf BUFF1_1149 (N3977, N3865_t1);
buf BUFF1_1150 (N3980, N3868_t0);
buf BUFF1_1151 (N3983, N3868_t1);
nand NAND2_1152 (N3987, N3924, N3925);
nand NAND4_1153 (N3992, N3765, N3894, N3930, N3931);
nand NAND4_1154 (N3996, N3766, N3895, N3935, N3936);
not NOT1_1155 (N4013, N3921_t0);
and AND2_1156 (N4028, N3932_t0, N3926_t0);
nand NAND2_1157 (N4029, N3953_t0, N3681);
nand NAND2_1158 (N4030, N3959_t0, N3686);
nand NAND2_1159 (N4031, N3965_t0, N3688);
nand NAND2_1160 (N4032, N3971_t0, N3689);
nand NAND2_1161 (N4033, N3977_t0, N3693);
nand NAND2_1162 (N4034, N3983_t0, N3695);
buf BUFF1_1163 (N4035, N3926_t1);
not NOT1_1164 (N4042, N3953_t1);
not NOT1_1165 (N4043, N3956_t0);
nand NAND2_1166 (N4044, N3956_t1, N3685);
not NOT1_1167 (N4045, N3959_t1);
not NOT1_1168 (N4046, N3962_t0);
nand NAND2_1169 (N4047, N3962_t1, N3687);
not NOT1_1170 (N4048, N3965_t1);
not NOT1_1171 (N4049, N3971_t1);
not NOT1_1172 (N4050, N3977_t1);
not NOT1_1173 (N4051, N3980_t0);
nand NAND2_1174 (N4052, N3980_t1, N3694);
not NOT1_1175 (N4053, N3983_t1);
not NOT1_1176 (N4054, N3974_t0);
nand NAND2_1177 (N4055, N3974_t1, N3696);
and AND2_1178 (N4056, N3932_t1, N2304_t1);
not NOT1_1179 (N4057, N3950_t0);
nand NAND2_1180 (N4058, N3950_t1, N3703);
buf BUFF1_1181 (N4059, N3937_t0);
buf BUFF1_1182 (N4062, N3937_t1);
not NOT1_1183 (N4065, N3968_t0);
nand NAND2_1184 (N4066, N3968_t1, N3704);
buf BUFF1_1185 (N4067, N3940_t0);
buf BUFF1_1186 (N4070, N3940_t1);
nand NAND2_1187 (N4073, N3926_t2, N3996_t0);
not NOT1_1188 (N4074, N3992_t0);
nand NAND2_1189 (N4075, N3493_t1, N4042);
nand NAND2_1190 (N4076, N3499_t1, N4045);
nand NAND2_1191 (N4077, N3505_t1, N4048);
nand NAND2_1192 (N4078, N3511_t1, N4049);
nand NAND2_1193 (N4079, N3517_t1, N4050);
nand NAND2_1194 (N4080, N3523_t1, N4053);
nand NAND2_1195 (N4085, N3496_t1, N4043);
nand NAND2_1196 (N4086, N3502_t1, N4046);
nand NAND2_1197 (N4088, N3520_t1, N4051);
nand NAND2_1198 (N4090, N3514_t1, N4054);
and AND2_1199 (N4091, N3996_t1, N1926_t2);
or OR2_1200 (N4094, N3605, N4056);
nand NAND2_1201 (N4098, N3490_t1, N4057);
nand NAND2_1202 (N4101, N3508_t1, N4065);
and AND2_1203 (N4104, N4073, N4074);
nand NAND2_1204 (N4105, N4075, N4029);
nand NAND2_1205 (N4106, N4062_t0, N3899);
nand NAND2_1206 (N4107, N4076, N4030);
nand NAND2_1207 (N4108, N4077, N4031);
nand NAND2_1208 (N4109, N4078, N4032);
nand NAND2_1209 (N4110, N4070_t0, N3906);
nand NAND2_1210 (N4111, N4079, N4033);
nand NAND2_1211 (N4112, N4080, N4034);
not NOT1_1212 (N4113, N4059_t0);
nand NAND2_1213 (N4114, N4059_t1, N3898);
not NOT1_1214 (N4115, N4062_t1);
nand NAND2_1215 (N4116, N4085, N4044);
nand NAND2_1216 (N4119, N4086, N4047);
not NOT1_1217 (N4122, N4070_t1);
nand NAND2_1218 (N4123, N4088, N4052);
not NOT1_1219 (N4126, N4067_t0);
nand NAND2_1220 (N4127, N4067_t1, N3911);
nand NAND2_1221 (N4128, N4090, N4055);
nand NAND2_1222 (N4139, N4098, N4058);
nand NAND2_1223 (N4142, N4101, N4066);
not NOT1_1224 (N4145, N4104);
not NOT1_1225 (N4146, N4105);
nand NAND2_1226 (N4147, N3824_t1, N4115);
not NOT1_1227 (N4148, N4107);
not NOT1_1228 (N4149, N4108);
not NOT1_1229 (N4150, N4109);
nand NAND2_1230 (N4151, N3830_t1, N4122);
not NOT1_1231 (N4152, N4111);
not NOT1_1232 (N4153, N4112);
nand NAND2_1233 (N4154, N3821_t1, N4113);
nand NAND2_1234 (N4161, N3827_t1, N4126);
buf BUFF1_1235 (N4167, N4091_t0);
buf BUFF1_1236 (N4174, N4094_t0);
buf BUFF1_1237 (N4182, N4091_t1);
and AND2_1238 (N4186, N330_t1, N4094_t1);
and AND2_1239 (N4189, N4146, N2230);
nand NAND2_1240 (N4190, N4147, N4106);
and AND2_1241 (N4191, N4148, N2232);
and AND2_1242 (N4192, N4149, N2233);
and AND2_1243 (N4193, N4150, N2234);
nand NAND2_1244 (N4194, N4151, N4110);
and AND2_1245 (N4195, N4152, N2236);
and AND2_1246 (N4196, N4153, N2237);
nand NAND2_1247 (N4197, N4154, N4114);
buf BUFF1_1248 (N4200, N4116_t0);
buf BUFF1_1249 (N4203, N4116_t1);
buf BUFF1_1250 (N4209, N4119_t0);
buf BUFF1_1251 (N4213, N4119_t1);
nand NAND2_1252 (N4218, N4161, N4127);
buf BUFF1_1253 (N4223, N4123_t0);
and AND2_1254 (N4238, N4128_t0, N3917_t0);
not NOT1_1255 (N4239, N4139_t0);
not NOT1_1256 (N4241, N4142_t0);
and AND2_1257 (N4242, N330_t2, N4123_t1);
buf BUFF1_1258 (N4247, N4128_t1);
nor NOR3_1259 (N4251, N3713, N4189, N2898);
not NOT1_1260 (N4252, N4190);
nor NOR3_1261 (N4253, N3715, N4191, N2900);
nor NOR3_1262 (N4254, N3716, N4192, N2901);
nor NOR3_1263 (N4255, N3717, N4193, N3406);
not NOT1_1264 (N4256, N4194);
nor NOR3_1265 (N4257, N3719, N4195, N3779);
nor NOR3_1266 (N4258, N3720, N4196, N3780);
and AND2_1267 (N4283, N4167_t0, N4035_t0);
and AND2_1268 (N4284, N4174_t0, N4035_t1);
or OR2_1269 (N4287, N3815_t0, N4238);
not NOT1_1270 (N4291, N4186_t0);
not NOT1_1271 (N4295, N4167_t1);
buf BUFF1_1272 (N4296, N4167_t2);
not NOT1_1273 (N4299, N4182_t0);
and AND2_1274 (N4303, N4252, N2231);
and AND2_1275 (N4304, N4256, N2235);
buf BUFF1_1276 (N4305, N4197_t0);
or OR2_1277 (N4310, N3992_t1, N4283);
and AND3_1278 (N4316, N4174_t1, N4213_t0, N4203_t0);
and AND2_1279 (N4317, N4174_t2, N4209_t0);
and AND3_1280 (N4318, N4223_t0, N4128_t2, N4218_t0);
and AND2_1281 (N4319, N4223_t1, N4128_t3);
and AND2_1282 (N4322, N4167_t3, N4209_t1);
nand NAND2_1283 (N4325, N4203_t1, N3913_t0);
nand NAND3_1284 (N4326, N4203_t2, N4213_t1, N4167_t4);
nand NAND2_1285 (N4327, N4218_t1, N3815_t1);
nand NAND3_1286 (N4328, N4218_t2, N4128_t4, N3917_t1);
nand NAND2_1287 (N4329, N4247_t0, N4013);
not NOT1_1288 (N4330, N4247_t1);
and AND3_1289 (N4331, N330_t3, N4094_t2, N4295);
and AND2_1290 (N4335, N4251, N2730);
and AND2_1291 (N4338, N4253, N2734);
and AND2_1292 (N4341, N4254, N2736);
and AND2_1293 (N4344, N4255, N2738);
and AND2_1294 (N4347, N4257, N2742);
and AND2_1295 (N4350, N4258, N2744);
buf BUFF1_1296 (N4353, N4197_t1);
buf BUFF1_1297 (N4356, N4203_t3);
buf BUFF1_1298 (N4359, N4209_t2);
buf BUFF1_1299 (N4362, N4218_t3);
buf BUFF1_1300 (N4365, N4242_t0);
buf BUFF1_1301 (N4368, N4242_t1);
and AND2_1302 (N4371, N4223_t2, N4223);
nor NOR3_1303 (N4376, N3714, N4303, N2899);
nor NOR3_1304 (N4377, N3718, N4304, N3642);
and AND2_1305 (N4387, N330_t4, N4317);
and AND2_1306 (N4390, N330_t5, N4318);
nand NAND2_1307 (N4393, N3921_t1, N4330);
buf BUFF1_1308 (N4398, N4287_t0);
buf BUFF1_1309 (N4413, N4284_t0);
nand NAND3_1310 (N4416, N3920, N4325, N4326);
or OR2_1311 (N4421, N3812_t1, N4322);
nand NAND3_1312 (N4427, N3948, N4327, N4328);
buf BUFF1_1313 (N4430, N4287_t1);
and AND2_1314 (N4435, N330_t6, N4316);
or OR2_1315 (N4442, N4331_t0, N4296_t0);
and AND4_1316 (N4443, N4174_t3, N4305_t0, N4203_t4, N4213_t2);
nand NAND2_1317 (N4446, N4305_t1, N3809_t1);
nand NAND3_1318 (N4447, N4305_t2, N4200_t0, N3913_t1);
nand NAND4_1319 (N4448, N4305_t3, N4200_t1, N4213_t3, N4167_t5);
not NOT1_1320 (N4452, N4356_t0);
nand NAND2_1321 (N4458, N4329, N4393);
not NOT1_1322 (N4461, N4365_t0);
not NOT1_1323 (N4462, N4368_t0);
nand NAND2_1324 (N4463, N4371_t0, N1460);
not NOT1_1325 (N4464, N4371_t1);
buf BUFF1_1326 (N4465, N4310_t0);
nor NOR2_1327 (N4468, N4331_t1, N4296_t1);
and AND2_1328 (N4472, N4376, N2732);
and AND2_1329 (N4475, N4377, N2740);
buf BUFF1_1330 (N4479, N4310_t1);
not NOT1_1331 (N4484, N4353_t0);
not NOT1_1332 (N4486, N4359_t0);
nand NAND2_1333 (N4487, N4359_t1, N4299);
not NOT1_1334 (N4491, N4362_t0);
and AND2_1335 (N4493, N330_t7, N4319_t0);
not NOT1_1336 (N4496, N4398_t0);
and AND2_1337 (N4497, N4287_t2, N4398_t1);
and AND2_1338 (N4498, N4442, N1769);
nand NAND4_1339 (N4503, N3947, N4446, N4447, N4448);
not NOT1_1340 (N4506, N4413_t0);
not NOT1_1341 (N4507, N4435_t0);
not NOT1_1342 (N4508, N4421_t0);
nand NAND2_1343 (N4509, N4421_t1, N4452);
not NOT1_1344 (N4510, N4427_t0);
nand NAND2_1345 (N4511, N4427_t1, N4241);
nand NAND2_1346 (N4515, N965_t1, N4464);
not NOT1_1347 (N4526, N4416_t0);
nand NAND2_1348 (N4527, N4416_t1, N4484);
nand NAND2_1349 (N4528, N4182_t1, N4486);
not NOT1_1350 (N4529, N4430_t0);
nand NAND2_1351 (N4530, N4430_t1, N4491);
buf BUFF1_1352 (N4531, N4387_t0);
buf BUFF1_1353 (N4534, N4387_t1);
buf BUFF1_1354 (N4537, N4390_t0);
buf BUFF1_1355 (N4540, N4390_t1);
and AND3_1356 (N4545, N330_t8, N4319_t1, N4496);
and AND2_1357 (N4549, N330_t9, N4443_t0);
nand NAND2_1358 (N4552, N4356_t1, N4508);
nand NAND2_1359 (N4555, N4142_t1, N4510);
not NOT1_1360 (N4558, N4493_t0);
nand NAND2_1361 (N4559, N4463, N4515);
not NOT1_1362 (N4562, N4465_t0);
and AND2_1363 (N4563, N4310_t2, N4465_t1);
buf BUFF1_1364 (N4564, N4468_t0);
not NOT1_1365 (N4568, N4479_t0);
buf BUFF1_1366 (N4569, N4443_t1);
nand NAND2_1367 (N4572, N4353_t1, N4526);
nand NAND2_1368 (N4573, N4362_t1, N4529);
nand NAND2_1369 (N4576, N4487, N4528);
buf BUFF1_1370 (N4581, N4458_t0);
buf BUFF1_1371 (N4584, N4458_t1);
or OR3_1372 (N4587, N2758_t0, N4498_t0, N2761_t0);
nor NOR3_1373 (N4588, N2758_t1, N4498_t1, N2761_t1);
or OR2_1374 (N4589, N4545, N4497);
nand NAND2_1375 (N4593, N4552, N4509);
not NOT1_1376 (N4596, N4531_t0);
not NOT1_1377 (N4597, N4534_t0);
nand NAND2_1378 (N4599, N4555, N4511);
not NOT1_1379 (N4602, N4537_t0);
not NOT1_1380 (N4603, N4540_t0);
and AND3_1381 (N4608, N330_t10, N4284_t1, N4562);
buf BUFF1_1382 (N4613, N4503_t0);
buf BUFF1_1383 (N4616, N4503_t1);
nand NAND2_1384 (N4619, N4572, N4527);
nand NAND2_1385 (N4623, N4573, N4530);
not NOT1_1386 (N4628, N4588);
nand NAND2_1387 (N4629, N4569_t0, N4506);
not NOT1_1388 (N4630, N4569_t1);
not NOT1_1389 (N4635, N4576_t0);
nand NAND2_1390 (N4636, N4576_t1, N4291);
not NOT1_1391 (N4640, N4581_t0);
nand NAND2_1392 (N4641, N4581_t1, N4461);
not NOT1_1393 (N4642, N4584_t0);
nand NAND2_1394 (N4643, N4584_t1, N4462);
nor NOR2_1395 (N4644, N4608, N4563);
and AND2_1396 (N4647, N4559_t0, N2128);
and AND2_1397 (N4650, N4559_t1, N2743);
buf BUFF1_1398 (N4656, N4549_t0);
buf BUFF1_1399 (N4659, N4549_t1);
buf BUFF1_1400 (N4664, N4564_t0);
and AND2_1401 (N4667, N4587, N4628);
nand NAND2_1402 (N4668, N4413_t1, N4630);
not NOT1_1403 (N4669, N4616_t0);
nand NAND2_1404 (N4670, N4616_t1, N4239);
not NOT1_1405 (N4673, N4619_t0);
nand NAND2_1406 (N4674, N4619_t1, N4507);
nand NAND2_1407 (N4675, N4186_t1, N4635);
not NOT1_1408 (N4676, N4623_t0);
nand NAND2_1409 (N4677, N4623_t1, N4558);
nand NAND2_1410 (N4678, N4365_t1, N4640);
nand NAND2_1411 (N4679, N4368_t1, N4642);
not NOT1_1412 (N4687, N4613_t0);
nand NAND2_1413 (N4688, N4613_t1, N4568);
buf BUFF1_1414 (N4691, N4593_t0);
buf BUFF1_1415 (N4694, N4593_t1);
buf BUFF1_1416 (N4697, N4599_t0);
buf BUFF1_1417 (N4700, N4599_t1);
nand NAND2_1418 (N4704, N4629, N4668);
nand NAND2_1419 (N4705, N4139_t1, N4669);
not NOT1_1420 (N4706, N4656_t0);
not NOT1_1421 (N4707, N4659_t0);
nand NAND2_1422 (N4708, N4435_t1, N4673);
nand NAND2_1423 (N4711, N4675, N4636);
nand NAND2_1424 (N4716, N4493_t1, N4676);
nand NAND2_1425 (N4717, N4678, N4641);
nand NAND2_1426 (N4721, N4679, N4643);
buf BUFF1_1427 (N4722, N4644_t0);
not NOT1_1428 (N4726, N4664_t0);
or OR3_1429 (N4727, N4647_t0, N4650_t0, N4350_t0);
nor NOR3_1430 (N4730, N4647_t1, N4650_t1, N4350_t1);
nand NAND2_1431 (N4733, N4479_t1, N4687);
nand NAND2_1432 (N4740, N4705, N4670);
nand NAND2_1433 (N4743, N4708, N4674);
not NOT1_1434 (N4747, N4691_t0);
nand NAND2_1435 (N4748, N4691_t1, N4596);
not NOT1_1436 (N4749, N4694_t0);
nand NAND2_1437 (N4750, N4694_t1, N4597);
not NOT1_1438 (N4753, N4697_t0);
nand NAND2_1439 (N4754, N4697_t1, N4602);
not NOT1_1440 (N4755, N4700_t0);
nand NAND2_1441 (N4756, N4700_t1, N4603);
nand NAND2_1442 (N4757, N4716, N4677);
nand NAND2_1443 (N4769, N4733, N4688);
and AND2_1444 (N4772, N330_t11, N4704);
not NOT1_1445 (N4775, N4721);
not NOT1_1446 (N4778, N4730_t0);
nand NAND2_1447 (N4786, N4531_t1, N4747);
nand NAND2_1448 (N4787, N4534_t1, N4749);
nand NAND2_1449 (N4788, N4537_t1, N4753);
nand NAND2_1450 (N4789, N4540_t1, N4755);
and AND2_1451 (N4794, N4711_t0, N2124);
and AND2_1452 (N4797, N4711_t1, N2735);
and AND2_1453 (N4800, N4717_t0, N2127);
buf BUFF1_1454 (N4805, N4722_t0);
and AND2_1455 (N4808, N4717_t1, N4468_t1);
buf BUFF1_1456 (N4812, N4727_t0);
and AND2_1457 (N4815, N4727_t1, N4778);
not NOT1_1458 (N4816, N4769_t0);
not NOT1_1459 (N4817, N4772_t0);
nand NAND2_1460 (N4818, N4786, N4748);
nand NAND2_1461 (N4822, N4787, N4750);
nand NAND2_1462 (N4823, N4788, N4754);
nand NAND2_1463 (N4826, N4789, N4756);
nand NAND2_1464 (N4829, N4775_t0, N4726);
not NOT1_1465 (N4830, N4775_t1);
and AND2_1466 (N4831, N4743_t0, N2122);
and AND2_1467 (N4838, N4757_t0, N2126);
buf BUFF1_1468 (N4844, N4740_t0);
buf BUFF1_1469 (N4847, N4740_t1);
buf BUFF1_1470 (N4850, N4743_t1);
buf BUFF1_1471 (N4854, N4757_t1);
nand NAND2_1472 (N4859, N4772_t1, N4816);
nand NAND2_1473 (N4860, N4769_t1, N4817);
not NOT1_1474 (N4868, N4826);
not NOT1_1475 (N4870, N4805_t0);
not NOT1_1476 (N4872, N4808_t0);
nand NAND2_1477 (N4873, N4664_t1, N4830);
or OR3_1478 (N4876, N4794_t0, N4797_t0, N4341_t0);
nor NOR3_1479 (N4880, N4794_t1, N4797_t1, N4341_t1);
not NOT1_1480 (N4885, N4812_t0);
not NOT1_1481 (N4889, N4822);
nand NAND2_1482 (N4895, N4859, N4860);
not NOT1_1483 (N4896, N4844_t0);
nand NAND2_1484 (N4897, N4844_t1, N4706);
not NOT1_1485 (N4898, N4847_t0);
nand NAND2_1486 (N4899, N4847_t1, N4707);
nor NOR2_1487 (N4900, N4868, N4564_t1);
and AND4_1488 (N4901, N4717_t2, N4757_t2, N4823_t0, N4564_t2);
not NOT1_1489 (N4902, N4850_t0);
not NOT1_1490 (N4904, N4854_t0);
nand NAND2_1491 (N4905, N4854_t1, N4872);
nand NAND2_1492 (N4906, N4873, N4829);
and AND2_1493 (N4907, N4818_t0, N2123);
and AND2_1494 (N4913, N4823_t1, N2125);
and AND2_1495 (N4916, N4818_t1, N4644_t1);
not NOT1_1496 (N4920, N4880_t0);
and AND2_1497 (N4921, N4895, N2184);
nand NAND2_1498 (N4924, N4656_t1, N4896);
nand NAND2_1499 (N4925, N4659_t1, N4898);
or OR2_1500 (N4926, N4900, N4901);
nand NAND2_1501 (N4928, N4889_t0, N4870);
not NOT1_1502 (N4929, N4889_t1);
nand NAND2_1503 (N4930, N4808_t1, N4904);
not NOT1_1504 (N4931, N4906);
buf BUFF1_1505 (N4937, N4876_t0);
buf BUFF1_1506 (N4940, N4876_t1);
and AND2_1507 (N4944, N4876_t2, N4920);
nand NAND2_1508 (N4946, N4924, N4897);
nand NAND2_1509 (N4949, N4925, N4899);
nand NAND2_1510 (N4950, N4916_t0, N4902);
not NOT1_1511 (N4951, N4916_t1);
nand NAND2_1512 (N4952, N4805_t1, N4929);
nand NAND2_1513 (N4953, N4930, N4905);
and AND2_1514 (N4954, N4926, N2737);
and AND2_1515 (N4957, N4931, N2741);
or OR3_1516 (N4964, N2764_t0, N2483_t0, N4921_t0);
nor NOR3_1517 (N4965, N2764_t1, N2483_t1, N4921_t1);
not NOT1_1518 (N4968, N4949);
nand NAND2_1519 (N4969, N4850_t1, N4951);
nand NAND2_1520 (N4970, N4952, N4928);
and AND2_1521 (N4973, N4953, N2739);
not NOT1_1522 (N4978, N4937_t0);
not NOT1_1523 (N4979, N4940_t0);
not NOT1_1524 (N4980, N4965);
nor NOR2_1525 (N4981, N4968, N4722_t1);
and AND4_1526 (N4982, N4818_t2, N4743_t2, N4946_t0, N4722_t2);
nand NAND2_1527 (N4983, N4950, N4969);
not NOT1_1528 (N4984, N4970);
and AND2_1529 (N4985, N4946_t1, N2121);
or OR3_1530 (N4988, N4913_t0, N4954_t0, N4344_t0);
nor NOR3_1531 (N4991, N4913_t1, N4954_t1, N4344_t1);
or OR3_1532 (N4996, N4800_t0, N4957_t0, N4347_t0);
nor NOR3_1533 (N4999, N4800_t1, N4957_t1, N4347_t1);
and AND2_1534 (N5002, N4964, N4980);
or OR2_1535 (N5007, N4981, N4982);
and AND2_1536 (N5010, N4983, N2731);
and AND2_1537 (N5013, N4984, N2733);
or OR3_1538 (N5018, N4838_t0, N4973_t0, N4475_t0);
nor NOR3_1539 (N5021, N4838_t1, N4973_t1, N4475_t1);
not NOT1_1540 (N5026, N4991_t0);
not NOT1_1541 (N5029, N4999_t0);
and AND2_1542 (N5030, N5007, N2729);
buf BUFF1_1543 (N5039, N4996_t0);
buf BUFF1_1544 (N5042, N4988_t0);
and AND2_1545 (N5045, N4988_t1, N5026);
not NOT1_1546 (N5046, N5021_t0);
and AND2_1547 (N5047, N4996_t1, N5029);
or OR3_1548 (N5050, N4831_t0, N5010_t0, N4472_t0);
nor NOR3_1549 (N5055, N4831_t1, N5010_t1, N4472_t1);
or OR3_1550 (N5058, N4907_t0, N5013_t0, N4338_t0);
nor NOR3_1551 (N5061, N4907_t1, N5013_t1, N4338_t1);
and AND4_1552 (N5066, N4730_t1, N4999_t1, N5021_t1, N4991_t1);
buf BUFF1_1553 (N5070, N5018_t0);
and AND2_1554 (N5078, N5018_t1, N5046);
or OR3_1555 (N5080, N4985_t0, N5030_t0, N4335_t0);
nor NOR3_1556 (N5085, N4985_t1, N5030_t1, N4335_t1);
nand NAND2_1557 (N5094, N5039_t0, N4885);
not NOT1_1558 (N5095, N5039_t1);
not NOT1_1559 (N5097, N5042_t0);
and AND2_1560 (N5102, N5050_t0, N5050);
not NOT1_1561 (N5103, N5061_t0);
nand NAND2_1562 (N5108, N4812_t1, N5095);
not NOT1_1563 (N5109, N5070_t0);
nand NAND2_1564 (N5110, N5070_t1, N5097);
buf BUFF1_1565 (N5111, N5058_t0);
and AND2_1566 (N5114, N5050_t1, N1461_t0);
buf BUFF1_1567 (N5117, N5050_t2);
and AND2_1568 (N5120, N5080_t0, N5080);
and AND2_1569 (N5121, N5058_t1, N5103);
nand NAND2_1570 (N5122, N5094, N5108);
nand NAND2_1571 (N5125, N5042_t1, N5109);
and AND2_1572 (N5128, N1461_t1, N5080_t1);
and AND4_1573 (N5133, N4880_t1, N5061_t1, N5055_t0, N5085_t0);
and AND3_1574 (N5136, N5055_t1, N5085_t1, N1464_t1);
buf BUFF1_1575 (N5139, N5080_t2);
nand NAND2_1576 (N5145, N5125, N5110);
buf BUFF1_1577 (N5151, N5111_t0);
buf BUFF1_1578 (N5154, N5111_t1);
not NOT1_1579 (N5159, N5117_t0);
buf BUFF1_1580 (N5160, N5114_t0);
buf BUFF1_1581 (N5163, N5114_t1);
and AND2_1582 (N5166, N5066_t0, N5133_t0);
and AND2_1583 (N5173, N5066_t1, N5133_t1);
buf BUFF1_1584 (N5174, N5122_t0);
buf BUFF1_1585 (N5177, N5122_t1);
not NOT1_1586 (N5182, N5139_t0);
nand NAND2_1587 (N5183, N5139_t1, N5159);
buf BUFF1_1588 (N5184, N5128_t0);
buf BUFF1_1589 (N5188, N5128_t1);
not NOT1_1590 (N5192, N5166);
nor NOR2_1591 (N5193, N5136, N5173);
nand NAND2_1592 (N5196, N5151_t0, N4978);
not NOT1_1593 (N5197, N5151_t1);
nand NAND2_1594 (N5198, N5154_t0, N4979);
not NOT1_1595 (N5199, N5154_t1);
not NOT1_1596 (N5201, N5160_t0);
not NOT1_1597 (N5203, N5163_t0);
buf BUFF1_1598 (N5205, N5145_t0);
buf BUFF1_1599 (N5209, N5145_t1);
nand NAND2_1600 (N5212, N5117_t1, N5182);
and AND2_1601 (N5215, N213_t7, N5193);
not NOT1_1602 (N5217, N5174_t0);
not NOT1_1603 (N5219, N5177_t0);
nand NAND2_1604 (N5220, N4937_t1, N5197);
nand NAND2_1605 (N5221, N4940_t1, N5199);
not NOT1_1606 (N5222, N5184_t0);
nand NAND2_1607 (N5223, N5184_t1, N5201);
nand NAND2_1608 (N5224, N5188_t0, N5203);
not NOT1_1609 (N5225, N5188_t1);
nand NAND2_1610 (N5228, N5183, N5212);
not NOT1_1611 (N5231, N5215);
nand NAND2_1612 (N5232, N5205_t0, N5217);
not NOT1_1613 (N5233, N5205_t1);
nand NAND2_1614 (N5234, N5209_t0, N5219);
not NOT1_1615 (N5235, N5209_t1);
nand NAND2_1616 (N5236, N5196, N5220);
nand NAND2_1617 (N5240, N5198, N5221);
nand NAND2_1618 (N5242, N5160_t1, N5222);
nand NAND2_1619 (N5243, N5163_t1, N5225);
nand NAND2_1620 (N5245, N5174_t1, N5233);
nand NAND2_1621 (N5246, N5177_t1, N5235);
not NOT1_1622 (N5250, N5240);
not NOT1_1623 (N5253, N5228_t0);
nand NAND2_1624 (N5254, N5242, N5223);
nand NAND2_1625 (N5257, N5243, N5224);
nand NAND2_1626 (N5258, N5232, N5245);
nand NAND2_1627 (N5261, N5234, N5246);
not NOT1_1628 (N5266, N5257);
buf BUFF1_1629 (N5269, N5236_t0);
and AND3_1630 (N5277, N5236_t1, N5254_t0, N2307_t0);
and AND3_1631 (N5278, N5250_t0, N5254_t1, N2310_t0);
not NOT1_1632 (N5279, N5261);
not NOT1_1633 (N5283, N5269_t0);
nand NAND2_1634 (N5284, N5269_t1, N5253);
and AND3_1635 (N5285, N5236_t2, N5266_t0, N2310_t1);
and AND3_1636 (N5286, N5250_t1, N5266_t1, N2307_t1);
buf BUFF1_1637 (N5289, N5258_t0);
buf BUFF1_1638 (N5292, N5258_t1);
nand NAND2_1639 (N5295, N5228_t1, N5283);
or OR4_1640 (N5298, N5277, N5285, N5278, N5286);
buf BUFF1_1641 (N5303, N5279_t0);
buf BUFF1_1642 (N5306, N5279_t1);
nand NAND2_1643 (N5309, N5295, N5284);
not NOT1_1644 (N5312, N5292_t0);
not NOT1_1645 (N5313, N5289_t0);
not NOT1_1646 (N5322, N5306_t0);
not NOT1_1647 (N5323, N5303_t0);
buf BUFF1_1648 (N5324, N5298_t0);
buf BUFF1_1649 (N5327, N5298_t1);
buf BUFF1_1650 (N5332, N5309_t0);
buf BUFF1_1651 (N5335, N5309_t1);
nand NAND2_1652 (N5340, N5324_t0, N5323);
nand NAND2_1653 (N5341, N5327_t0, N5322);
not NOT1_1654 (N5344, N5327_t1);
not NOT1_1655 (N5345, N5324_t1);
nand NAND2_1656 (N5348, N5332_t0, N5313);
nand NAND2_1657 (N5349, N5335_t0, N5312);
nand NAND2_1658 (N5350, N5303_t1, N5345);
nand NAND2_1659 (N5351, N5306_t1, N5344);
not NOT1_1660 (N5352, N5335_t1);
not NOT1_1661 (N5353, N5332_t1);
nand NAND2_1662 (N5354, N5289_t1, N5353);
nand NAND2_1663 (N5355, N5292_t1, N5352);
nand NAND2_1664 (N5356, N5350, N5340);
nand NAND2_1665 (N5357, N5351, N5341);
nand NAND2_1666 (N5358, N5348, N5354);
nand NAND2_1667 (N5359, N5349, N5355);
and AND2_1668 (N5360, N5356, N5357);
nand NAND2_1669 (N5361, N5358, N5359);

endmodule
