// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module c1908f (INC,END,clk,rst,N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;

output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N1_t0,N1_t1,N4_t0,N4_t1,N7_t0,N7_t1,N10_t0,N10_t1,N13_t0,
     N13_t1,N16_t0,N16_t1,N19_t0,N19_t1,N22_t0,N22_t1,N25_t0,N25_t1,N28_t0,
     N28_t1,N31_t0,N31_t1,N34_t0,N34_t1,N37_t0,N37_t1,N40_t0,N40_t1,N43_t0,
     N43_t1,N46_t0,N46_t1,N63_t0,N63_t1,N88_t0,N88_t1,N66_t0,N66_t1,N91_t0,
     N91_t1,N72_t0,N72_t1,N72_t2,N69_t0,N69_t1,N76_t0,N76_t1,N79_t0,N79_t1,
     N82_t0,N82_t1,N85_t0,N85_t1,N104_t0,N104_t1,N104_t2,N104_t3,N104_t4,N104_t5,
     N104_t6,N94_t0,N94_t1,N94_t2,N94_t3,N99_t0,N99_t1,N99_t2,N99_t3,N343_t0,
     N343_t1,N346_t0,N346_t1,N349_t0,N349_t1,N352_t0,N352_t1,N355_t0,N355_t1,N358_t0,
     N358_t1,N361_t0,N361_t1,N364_t0,N364_t1,N367_t0,N367_t1,N370_t0,N370_t1,N373_t0,
     N373_t1,N376_t0,N376_t1,N379_t0,N379_t1,N382_t0,N382_t1,N385_t0,N385_t1,N388_t0,
     N388_t1,N306_t0,N306_t1,N306_t2,N306_t3,N306_t4,N306_t5,N331_t0,N331_t1,N331_t2,
     N331_t3,N331_t4,N331_t5,N190_t0,N190_t1,N190_t2,N194_t0,N194_t1,N206_t0,N206_t1,
     N209_t0,N209_t1,N225_t0,N225_t1,N225_t2,N243_t0,N243_t1,N243_t2,N319_t0,N319_t1,
     N319_t2,N319_t3,N319_t4,N319_t5,N220_t0,N220_t1,N220_t2,N220_t3,N229_t0,N229_t1,
     N232_t0,N232_t1,N239_t0,N239_t1,N239_t2,N49_t0,N49_t1,N49_t2,N253_t0,N253_t1,
     N247_t0,N247_t1,N247_t2,N326_t0,N326_t1,N326_t2,N326_t3,N277_t0,N277_t1,N280_t0,
     N280_t1,N260_t0,N260_t1,N300_t0,N300_t1,N201_t0,N201_t1,N201_t2,N201_t3,N216_t0,
     N216_t1,N216_t2,N197_t0,N197_t1,N197_t2,N56_t0,N56_t1,N56_t2,N257_t0,N257_t1,
     N235_t0,N235_t1,N235_t2,N60_t0,N60_t1,N263_t0,N263_t1,N266_t0,N266_t1,N269_t0,
     N269_t1,N272_t0,N272_t1,N316_t0,N316_t1,N212_t0,N212_t1,N212_t2,N53_t0,N53_t1,
     N682_t0,N682_t1,N685_t0,N685_t1,N616_t0,N616_t1,N619_t0,N619_t1,N622_t0,N622_t1,
     N625_t0,N625_t1,N631_t0,N631_t1,N643_t0,N643_t1,N649_t0,N649_t1,N652_t0,N652_t1,
     N655_t0,N655_t1,N612_t0,N612_t1,N612_t2,N608_t0,N608_t1,N608_t2,N661_t0,N661_t1,
     N658_t0,N658_t1,N667_t0,N667_t1,N664_t0,N664_t1,N673_t0,N673_t1,N670_t0,N670_t1,
     N679_t0,N679_t1,N676_t0,N676_t1,N297_t0,N297_t1,N603_t0,N603_t1,N603_t2,N603_t3,
     N303_t0,N303_t1,N338_t0,N338_t1,N338_t2,N338_t3,N556_t0,N556_t1,N688_t0,N688_t1,
     N691_t0,N691_t1,N562_t0,N562_t1,N694_t0,N694_t1,N697_t0,N697_t1,N568_t0,N568_t1,
     N700_t0,N700_t1,N703_t0,N703_t1,N574_t0,N574_t1,N580_t0,N580_t1,N706_t0,N706_t1,
     N709_t0,N709_t1,N586_t0,N586_t1,N712_t0,N712_t1,N715_t0,N715_t1,N592_t0,N592_t1,
     N628_t0,N628_t1,N718_t0,N718_t1,N721_t0,N721_t1,N634_t0,N634_t1,N724_t0,N724_t1,
     N727_t0,N727_t1,N637_t0,N637_t1,N595_t0,N595_t1,N730_t0,N730_t1,N733_t0,N733_t1,
     N736_t0,N736_t1,N739_t0,N739_t1,N640_t0,N640_t1,N742_t0,N742_t1,N745_t0,N745_t1,
     N646_t0,N646_t1,N748_t0,N748_t1,N751_t0,N751_t1,N559_t0,N559_t1,N565_t0,N565_t1,
     N571_t0,N571_t1,N577_t0,N577_t1,N583_t0,N583_t1,N589_t0,N589_t1,N598_t0,N598_t1,
     N939_t0,N939_t1,N935_t0,N935_t1,N943_t0,N943_t1,N947_t0,N947_t1,N955_t0,N955_t1,
     N951_t0,N951_t1,N962_t0,N962_t1,N969_t0,N969_t1,N977_t0,N977_t1,N985_t0,N985_t1,
     N998_t0,N998_t1,N899_t0,N899_t1,N899_t2,N903_t0,N903_t1,N903_t2,N923_t0,N923_t1,
     N1010_t0,N1010_t1,N1013_t0,N1013_t1,N1016_t0,N1016_t1,N1019_t0,N1019_t1,N1022_t0,N1022_t1,
     N1025_t0,N1025_t1,N1028_t0,N1028_t1,N959_t0,N959_t1,N1031_t0,N1031_t1,N1034_t0,N1034_t1,
     N965_t0,N965_t1,N1037_t0,N1037_t1,N1040_t0,N1040_t1,N973_t0,N973_t1,N1043_t0,N1043_t1,
     N981_t0,N981_t1,N1046_t0,N1046_t1,N994_t0,N994_t1,N1049_t0,N1049_t1,N907_t0,N907_t1,
     N910_t0,N910_t1,N1249_t0,N1249_t1,N1255_t0,N1255_t1,N1252_t0,N1252_t1,N1261_t0,N1261_t1,
     N1258_t0,N1258_t1,N1232_t0,N1232_t1,N1235_t0,N1235_t1,N1243_t0,N1243_t1,N1246_t0,N1246_t1,
     N1319_t0,N1319_t1,N1334_t0,N1334_t1,N1264_t0,N1264_t1,N1355_t0,N1355_t1,N1352_t0,N1352_t1,
     N1358_t0,N1358_t1,N1361_t0,N1361_t1,N1367_t0,N1367_t1,N1364_t0,N1364_t1,N1373_t0,N1373_t1,
     N1379_t0,N1379_t1,N1383_t0,N1383_t1,N1393_t0,N1393_t1,N1370_t0,N1370_t1,N1376_t0,N1376_t1,
     N1390_t0,N1390_t1,N1419_t0,N1419_t1,N1416_t0,N1416_t1,N1440_t0,N1440_t1,N1472_t0,N1472_t1,
     N1478_t0,N1478_t1,N1481_t0,N1481_t1,N1484_t0,N1484_t1,N1510_t0,N1510_t1,N1522_t0,N1522_t1,
     N1522_t2,N1534_t0,N1534_t1,N1537_t0,N1537_t1,N1540_t0,N1540_t1,N1517_t0,N1517_t1,N1514_t0,
     N1514_t1,N1557_t0,N1557_t1,N1557_t2,N1554_t0,N1554_t1,N1571_t0,N1571_t1,N1576_t0,N1576_t1,
     N1561_t0,N1561_t1,N1546_t0,N1546_t1,N1596_t0,N1596_t1,N1600_t0,N1600_t1,N1603_t0,N1603_t1,
     N1606_t0,N1606_t1,N1609_t0,N1609_t1,N1612_t0,N1612_t1,N1615_t0,N1615_t1,N1588_t0,N1588_t1,
     N1643_t0,N1643_t1,N1647_t0,N1647_t1,N1651_t0,N1651_t1,N1620_t0,N1620_t1,N1658_t0,N1658_t1,
     N1661_t0,N1661_t1,N1640_t0,N1640_t1,N1664_t0,N1664_t1,N1623_t0,N1623_t1,N1685_t0,N1685_t1,
     N1697_t0,N1697_t1,N1701_t0,N1701_t1,N1717_t0,N1717_t1,N1723_t0,N1723_t1,N1731_t0,N1731_t1,
     N1714_t0,N1714_t1,N1734_t0,N1734_t1,N1751_t0,N1751_t1,N1742_t0,N1742_t1,N290_t0,N290_t1,
     N290_t2,N290_t3,N290_t4,N290_t5,N1748_t0,N1748_t1,N1777_t0,N1777_t1,N1774_t0,N1774_t1,
     N1788_t0,N1788_t1,N1815_t0,N1815_t1,N1818_t0,N1818_t1,N1798_t0,N1798_t1,N1812_t0,N1812_t1,
     N1802_t0,N1802_t1,N1841_t0,N1841_t1,N1830_t0,N1830_t1,N1838_t0,N1838_t1,N1866_t0,N1866_t1,
     N1872_t0,N1872_t1,N1869_t0,N1869_t1,N1875_t0,N1875_t1,N1858_t0,N1858_t1,N1898_t0,N1898_t1,
     N1902_t0,N1902_t1,N1879_t0,N1879_t1,N1889_t0,N1889_t1,N1930_t0,N1930_t1,N1927_t0,N1927_t1,
     N1933_t0,N1933_t1,N1944_t0,N1944_t1,N1947_t0,N1947_t1,N1953_t0,N1953_t1,N1950_t0,N1950_t1,
     N1958_t0,N1958_t1,N1961_t0,N1961_t1,N1965_t0,N1965_t1,N1968_t0,N1968_t1,N1987_t0,N1987_t1,
     N1980_t0,N1980_t1,N2027_t0,N2027_t1,N2052_t0,N2052_t1,N2055_t0,N2055_t1,N2042_t0,N2042_t1,
     N2030_t0,N2030_t1,N2068_t0,N2068_t1,N2033_t0,N2033_t1,N2071_t0,N2071_t1,N2062_t0,N2062_t1,
     N2078_t0,N2078_t1,N2081_t0,N2081_t1,N2151_t0,N2151_t1,N2148_t0,N2148_t1,N2199_t0,N2199_t1,
     N2196_t0,N2196_t1,N2205_t0,N2205_t1,N2202_t0,N2202_t1,N2237_t0,N2237_t1,N2241_t0,N2241_t1,
     N1164_t0,N1164_t1,N2245_t0,N2245_t1,N1168_t0,N1168_t1,N2266_t0,N2266_t1,N2272_t0,N2272_t1,
     N2086_t0,N2086_t1,N2257_t0,N2257_t1,N2089_t0,N2089_t1,N2260_t0,N2260_t1,N2279_t0,N2279_t1,
     N313_t0,N313_t1,N2263_t0,N2263_t1,N2269_t0,N2269_t1,N2286_t0,N2286_t1,N2286_t2,N2286_t3,
     N2286_t4,N2286_t5,N2286_t6,N2286_t7,N2286_t8,N2286_t9,N2315_t0,N2315_t1,N2315_t2,N2315_t3,
     N2315_t4,N2315_t5,N2315_t6,N2315_t7,N2315_t8,N2315_t9,N2361_t0,N2361_t1,N2361_t2,N2361_t3,
     N2361_t4,N2361_t5,N2361_t6,N2361_t7,N2361_t8,N2361_t9,N2361_t10,N2361_t11,N2361_t12,N2104_t0,
     N2104_t1,N2104_t2,N2104_t3,N2104_t4,N2104_t5,N2104_t6,N2104_t7,N2104_t8,N2104_t9,N2104_t10,
     N2104_t11,N2104_t12,N2104_t13,N1171_t0,N1171_t1,N1171_t2,N1171_t3,N1171_t4,N1171_t5,N1171_t6,
     N1171_t7,N1171_t8,N1171_t9,N1171_t10,N1171_t11,N1171_t12,N1171_t13,N1171_t14,N1171_t15,N2340_t0,
     N2340_t1,N2340_t2,N2340_t3,N2340_t4,N2340_t5,N2340_t6,N2340_t7,N2340_t8,N2340_t9,N2340_t10,
     N2340_t11,N2129_t0,N2129_t1,N2129_t2,N2129_t3,N2129_t4,N2129_t5,N2129_t6,N2129_t7,N2129_t8,
     N2129_t9,N2129_t10,N2129_t11,N2129_t12,N2119_t0,N2119_t1,N2119_t2,N2119_t3,N2119_t4,N2119_t5,
     N2119_t6,N2119_t7,N2119_t8,N2353_t0,N2353_t1,N2353_t2,N2353_t3,N2353_t4,N2353_t5,N2353_t6,
     N2297_t0,N2297_t1,N2297_t2,N2297_t3,N2297_t4,N2297_t5,N2297_t6,N2297_t7,N2297_t8,N2297_t9,
     N2297_t10,N2297_t11,N2297_t12,N2297_t13,N2297_t14,N2375_t0,N2375_t1,N2375_t2,N2375_t3,N2375_t4,
     N2375_t5,N2375_t6,N2375_t7,N1188_t0,N1188_t1,N1188_t2,N1188_t3,N1188_t4,N1188_t5,N1188_t6,
     N1188_t7,N1188_t8,N1188_t9,N1188_t10,N1188_t11,N1188_t12,N1188_t13,N1188_t14,N1188_t15,N2326_t0,
     N2326_t1,N2326_t2,N2326_t3,N2326_t4,N2326_t5,N2326_t6,N2326_t7,N2326_t8,N2326_t9,N2326_t10,
     N2326_t11,N2326_t12,N2143_t0,N2143_t1,N2143_t2,N2143_t3,N2427_t0,N2427_t1,N2427_t2,N2427_t3,
     N2427_t4,N2427_t5,N2427_t6,N2427_t7,N2427_t8,N2427_t9,N2427_t10,N2427_t11,N2427_t12,N2427_t13,
     N2427_t14,N2427_t15,N2386_t0,N2386_t1,N2386_t2,N2386_t3,N2386_t4,N2386_t5,N2386_t6,N2386_t7,
     N2386_t8,N2386_t9,N2386_t10,N2386_t11,N2386_t12,N2386_t13,N926_t0,N926_t1,N926_t2,N926_t3,
     N926_t4,N926_t5,N926_t6,N926_t7,N2558_t0,N2558_t1,N2561_t0,N2561_t1,N2564_t0,N2564_t1,
     N2567_t0,N2567_t1,N2570_t0,N2570_t1,N2573_t0,N2573_t1,N2576_t0,N2576_t1,N2639_t0,N2639_t1,
     N2642_t0,N2642_t1,N2645_t0,N2645_t1,N2648_t0,N2648_t1,N2651_t0,N2651_t1,N2655_t0,N2655_t1,
     N2658_t0,N2658_t1,N2661_t0,N2661_t1,N2664_t0,N2664_t1,N2537_t0,N2537_t1,N2540_t0,N2540_t1,
     N2543_t0,N2543_t1,N2546_t0,N2546_t1,N2594_t0,N2594_t1,N2597_t0,N2597_t1,N2600_t0,N2600_t1,
     N2603_t0,N2603_t1,N2606_t0,N2606_t1,N2549_t0,N2549_t1,N2611_t0,N2611_t1,N2614_t0,N2614_t1,
     N2617_t0,N2617_t1,N2620_t0,N2620_t1,N2552_t0,N2552_t1,N2555_t0,N2555_t1,N2747_t0,N2747_t1,
     N2750_t0,N2750_t1,N2773_t0,N2773_t1,N2776_t0,N2776_t1,N283_t0,N283_t1,N283_t2,N283_t3,
     N283_t4,N283_t5,N2789_t0,N2789_t1,N2789_t2,N2789_t3,N2789_t4,N2789_t5,N2812_t0,N2812_t1,
     N2815_t0,N2815_t1,N2818_t0,N2818_t1,N2821_t0,N2821_t1,N2824_t0,N2824_t1,N2829_t0,N2829_t1,
     N2843_t0,N2843_t1,N2846_t0,N2846_t1,N2883_t0,N2883_t1;
reg [994:0] FEN;
fim FAN_N1_0 ( .fault(fault), .net(N1), .FEN(FEN[0]), .op(N1_t0) );
fim FAN_N1_1 ( .fault(fault), .net(N1), .FEN(FEN[1]), .op(N1_t1) );
fim FAN_N4_0 ( .fault(fault), .net(N4), .FEN(FEN[2]), .op(N4_t0) );
fim FAN_N4_1 ( .fault(fault), .net(N4), .FEN(FEN[3]), .op(N4_t1) );
fim FAN_N7_0 ( .fault(fault), .net(N7), .FEN(FEN[4]), .op(N7_t0) );
fim FAN_N7_1 ( .fault(fault), .net(N7), .FEN(FEN[5]), .op(N7_t1) );
fim FAN_N10_0 ( .fault(fault), .net(N10), .FEN(FEN[6]), .op(N10_t0) );
fim FAN_N10_1 ( .fault(fault), .net(N10), .FEN(FEN[7]), .op(N10_t1) );
fim FAN_N13_0 ( .fault(fault), .net(N13), .FEN(FEN[8]), .op(N13_t0) );
fim FAN_N13_1 ( .fault(fault), .net(N13), .FEN(FEN[9]), .op(N13_t1) );
fim FAN_N16_0 ( .fault(fault), .net(N16), .FEN(FEN[10]), .op(N16_t0) );
fim FAN_N16_1 ( .fault(fault), .net(N16), .FEN(FEN[11]), .op(N16_t1) );
fim FAN_N19_0 ( .fault(fault), .net(N19), .FEN(FEN[12]), .op(N19_t0) );
fim FAN_N19_1 ( .fault(fault), .net(N19), .FEN(FEN[13]), .op(N19_t1) );
fim FAN_N22_0 ( .fault(fault), .net(N22), .FEN(FEN[14]), .op(N22_t0) );
fim FAN_N22_1 ( .fault(fault), .net(N22), .FEN(FEN[15]), .op(N22_t1) );
fim FAN_N25_0 ( .fault(fault), .net(N25), .FEN(FEN[16]), .op(N25_t0) );
fim FAN_N25_1 ( .fault(fault), .net(N25), .FEN(FEN[17]), .op(N25_t1) );
fim FAN_N28_0 ( .fault(fault), .net(N28), .FEN(FEN[18]), .op(N28_t0) );
fim FAN_N28_1 ( .fault(fault), .net(N28), .FEN(FEN[19]), .op(N28_t1) );
fim FAN_N31_0 ( .fault(fault), .net(N31), .FEN(FEN[20]), .op(N31_t0) );
fim FAN_N31_1 ( .fault(fault), .net(N31), .FEN(FEN[21]), .op(N31_t1) );
fim FAN_N34_0 ( .fault(fault), .net(N34), .FEN(FEN[22]), .op(N34_t0) );
fim FAN_N34_1 ( .fault(fault), .net(N34), .FEN(FEN[23]), .op(N34_t1) );
fim FAN_N37_0 ( .fault(fault), .net(N37), .FEN(FEN[24]), .op(N37_t0) );
fim FAN_N37_1 ( .fault(fault), .net(N37), .FEN(FEN[25]), .op(N37_t1) );
fim FAN_N40_0 ( .fault(fault), .net(N40), .FEN(FEN[26]), .op(N40_t0) );
fim FAN_N40_1 ( .fault(fault), .net(N40), .FEN(FEN[27]), .op(N40_t1) );
fim FAN_N43_0 ( .fault(fault), .net(N43), .FEN(FEN[28]), .op(N43_t0) );
fim FAN_N43_1 ( .fault(fault), .net(N43), .FEN(FEN[29]), .op(N43_t1) );
fim FAN_N46_0 ( .fault(fault), .net(N46), .FEN(FEN[30]), .op(N46_t0) );
fim FAN_N46_1 ( .fault(fault), .net(N46), .FEN(FEN[31]), .op(N46_t1) );
fim FAN_N63_0 ( .fault(fault), .net(N63), .FEN(FEN[32]), .op(N63_t0) );
fim FAN_N63_1 ( .fault(fault), .net(N63), .FEN(FEN[33]), .op(N63_t1) );
fim FAN_N88_0 ( .fault(fault), .net(N88), .FEN(FEN[34]), .op(N88_t0) );
fim FAN_N88_1 ( .fault(fault), .net(N88), .FEN(FEN[35]), .op(N88_t1) );
fim FAN_N66_0 ( .fault(fault), .net(N66), .FEN(FEN[36]), .op(N66_t0) );
fim FAN_N66_1 ( .fault(fault), .net(N66), .FEN(FEN[37]), .op(N66_t1) );
fim FAN_N91_0 ( .fault(fault), .net(N91), .FEN(FEN[38]), .op(N91_t0) );
fim FAN_N91_1 ( .fault(fault), .net(N91), .FEN(FEN[39]), .op(N91_t1) );
fim FAN_N72_0 ( .fault(fault), .net(N72), .FEN(FEN[40]), .op(N72_t0) );
fim FAN_N72_1 ( .fault(fault), .net(N72), .FEN(FEN[41]), .op(N72_t1) );
fim FAN_N72_2 ( .fault(fault), .net(N72), .FEN(FEN[42]), .op(N72_t2) );
fim FAN_N69_0 ( .fault(fault), .net(N69), .FEN(FEN[43]), .op(N69_t0) );
fim FAN_N69_1 ( .fault(fault), .net(N69), .FEN(FEN[44]), .op(N69_t1) );
fim FAN_N76_0 ( .fault(fault), .net(N76), .FEN(FEN[45]), .op(N76_t0) );
fim FAN_N76_1 ( .fault(fault), .net(N76), .FEN(FEN[46]), .op(N76_t1) );
fim FAN_N79_0 ( .fault(fault), .net(N79), .FEN(FEN[47]), .op(N79_t0) );
fim FAN_N79_1 ( .fault(fault), .net(N79), .FEN(FEN[48]), .op(N79_t1) );
fim FAN_N82_0 ( .fault(fault), .net(N82), .FEN(FEN[49]), .op(N82_t0) );
fim FAN_N82_1 ( .fault(fault), .net(N82), .FEN(FEN[50]), .op(N82_t1) );
fim FAN_N85_0 ( .fault(fault), .net(N85), .FEN(FEN[51]), .op(N85_t0) );
fim FAN_N85_1 ( .fault(fault), .net(N85), .FEN(FEN[52]), .op(N85_t1) );
fim FAN_N104_0 ( .fault(fault), .net(N104), .FEN(FEN[53]), .op(N104_t0) );
fim FAN_N104_1 ( .fault(fault), .net(N104), .FEN(FEN[54]), .op(N104_t1) );
fim FAN_N104_2 ( .fault(fault), .net(N104), .FEN(FEN[55]), .op(N104_t2) );
fim FAN_N104_3 ( .fault(fault), .net(N104), .FEN(FEN[56]), .op(N104_t3) );
fim FAN_N104_4 ( .fault(fault), .net(N104), .FEN(FEN[57]), .op(N104_t4) );
fim FAN_N104_5 ( .fault(fault), .net(N104), .FEN(FEN[58]), .op(N104_t5) );
fim FAN_N104_6 ( .fault(fault), .net(N104), .FEN(FEN[59]), .op(N104_t6) );
fim FAN_N94_0 ( .fault(fault), .net(N94), .FEN(FEN[60]), .op(N94_t0) );
fim FAN_N94_1 ( .fault(fault), .net(N94), .FEN(FEN[61]), .op(N94_t1) );
fim FAN_N94_2 ( .fault(fault), .net(N94), .FEN(FEN[62]), .op(N94_t2) );
fim FAN_N94_3 ( .fault(fault), .net(N94), .FEN(FEN[63]), .op(N94_t3) );
fim FAN_N99_0 ( .fault(fault), .net(N99), .FEN(FEN[64]), .op(N99_t0) );
fim FAN_N99_1 ( .fault(fault), .net(N99), .FEN(FEN[65]), .op(N99_t1) );
fim FAN_N99_2 ( .fault(fault), .net(N99), .FEN(FEN[66]), .op(N99_t2) );
fim FAN_N99_3 ( .fault(fault), .net(N99), .FEN(FEN[67]), .op(N99_t3) );
fim FAN_N343_0 ( .fault(fault), .net(N343), .FEN(FEN[68]), .op(N343_t0) );
fim FAN_N343_1 ( .fault(fault), .net(N343), .FEN(FEN[69]), .op(N343_t1) );
fim FAN_N346_0 ( .fault(fault), .net(N346), .FEN(FEN[70]), .op(N346_t0) );
fim FAN_N346_1 ( .fault(fault), .net(N346), .FEN(FEN[71]), .op(N346_t1) );
fim FAN_N349_0 ( .fault(fault), .net(N349), .FEN(FEN[72]), .op(N349_t0) );
fim FAN_N349_1 ( .fault(fault), .net(N349), .FEN(FEN[73]), .op(N349_t1) );
fim FAN_N352_0 ( .fault(fault), .net(N352), .FEN(FEN[74]), .op(N352_t0) );
fim FAN_N352_1 ( .fault(fault), .net(N352), .FEN(FEN[75]), .op(N352_t1) );
fim FAN_N355_0 ( .fault(fault), .net(N355), .FEN(FEN[76]), .op(N355_t0) );
fim FAN_N355_1 ( .fault(fault), .net(N355), .FEN(FEN[77]), .op(N355_t1) );
fim FAN_N358_0 ( .fault(fault), .net(N358), .FEN(FEN[78]), .op(N358_t0) );
fim FAN_N358_1 ( .fault(fault), .net(N358), .FEN(FEN[79]), .op(N358_t1) );
fim FAN_N361_0 ( .fault(fault), .net(N361), .FEN(FEN[80]), .op(N361_t0) );
fim FAN_N361_1 ( .fault(fault), .net(N361), .FEN(FEN[81]), .op(N361_t1) );
fim FAN_N364_0 ( .fault(fault), .net(N364), .FEN(FEN[82]), .op(N364_t0) );
fim FAN_N364_1 ( .fault(fault), .net(N364), .FEN(FEN[83]), .op(N364_t1) );
fim FAN_N367_0 ( .fault(fault), .net(N367), .FEN(FEN[84]), .op(N367_t0) );
fim FAN_N367_1 ( .fault(fault), .net(N367), .FEN(FEN[85]), .op(N367_t1) );
fim FAN_N370_0 ( .fault(fault), .net(N370), .FEN(FEN[86]), .op(N370_t0) );
fim FAN_N370_1 ( .fault(fault), .net(N370), .FEN(FEN[87]), .op(N370_t1) );
fim FAN_N373_0 ( .fault(fault), .net(N373), .FEN(FEN[88]), .op(N373_t0) );
fim FAN_N373_1 ( .fault(fault), .net(N373), .FEN(FEN[89]), .op(N373_t1) );
fim FAN_N376_0 ( .fault(fault), .net(N376), .FEN(FEN[90]), .op(N376_t0) );
fim FAN_N376_1 ( .fault(fault), .net(N376), .FEN(FEN[91]), .op(N376_t1) );
fim FAN_N379_0 ( .fault(fault), .net(N379), .FEN(FEN[92]), .op(N379_t0) );
fim FAN_N379_1 ( .fault(fault), .net(N379), .FEN(FEN[93]), .op(N379_t1) );
fim FAN_N382_0 ( .fault(fault), .net(N382), .FEN(FEN[94]), .op(N382_t0) );
fim FAN_N382_1 ( .fault(fault), .net(N382), .FEN(FEN[95]), .op(N382_t1) );
fim FAN_N385_0 ( .fault(fault), .net(N385), .FEN(FEN[96]), .op(N385_t0) );
fim FAN_N385_1 ( .fault(fault), .net(N385), .FEN(FEN[97]), .op(N385_t1) );
fim FAN_N388_0 ( .fault(fault), .net(N388), .FEN(FEN[98]), .op(N388_t0) );
fim FAN_N388_1 ( .fault(fault), .net(N388), .FEN(FEN[99]), .op(N388_t1) );
fim FAN_N306_0 ( .fault(fault), .net(N306), .FEN(FEN[100]), .op(N306_t0) );
fim FAN_N306_1 ( .fault(fault), .net(N306), .FEN(FEN[101]), .op(N306_t1) );
fim FAN_N306_2 ( .fault(fault), .net(N306), .FEN(FEN[102]), .op(N306_t2) );
fim FAN_N306_3 ( .fault(fault), .net(N306), .FEN(FEN[103]), .op(N306_t3) );
fim FAN_N306_4 ( .fault(fault), .net(N306), .FEN(FEN[104]), .op(N306_t4) );
fim FAN_N306_5 ( .fault(fault), .net(N306), .FEN(FEN[105]), .op(N306_t5) );
fim FAN_N331_0 ( .fault(fault), .net(N331), .FEN(FEN[106]), .op(N331_t0) );
fim FAN_N331_1 ( .fault(fault), .net(N331), .FEN(FEN[107]), .op(N331_t1) );
fim FAN_N331_2 ( .fault(fault), .net(N331), .FEN(FEN[108]), .op(N331_t2) );
fim FAN_N331_3 ( .fault(fault), .net(N331), .FEN(FEN[109]), .op(N331_t3) );
fim FAN_N331_4 ( .fault(fault), .net(N331), .FEN(FEN[110]), .op(N331_t4) );
fim FAN_N331_5 ( .fault(fault), .net(N331), .FEN(FEN[111]), .op(N331_t5) );
fim FAN_N190_0 ( .fault(fault), .net(N190), .FEN(FEN[112]), .op(N190_t0) );
fim FAN_N190_1 ( .fault(fault), .net(N190), .FEN(FEN[113]), .op(N190_t1) );
fim FAN_N190_2 ( .fault(fault), .net(N190), .FEN(FEN[114]), .op(N190_t2) );
fim FAN_N194_0 ( .fault(fault), .net(N194), .FEN(FEN[115]), .op(N194_t0) );
fim FAN_N194_1 ( .fault(fault), .net(N194), .FEN(FEN[116]), .op(N194_t1) );
fim FAN_N206_0 ( .fault(fault), .net(N206), .FEN(FEN[117]), .op(N206_t0) );
fim FAN_N206_1 ( .fault(fault), .net(N206), .FEN(FEN[118]), .op(N206_t1) );
fim FAN_N209_0 ( .fault(fault), .net(N209), .FEN(FEN[119]), .op(N209_t0) );
fim FAN_N209_1 ( .fault(fault), .net(N209), .FEN(FEN[120]), .op(N209_t1) );
fim FAN_N225_0 ( .fault(fault), .net(N225), .FEN(FEN[121]), .op(N225_t0) );
fim FAN_N225_1 ( .fault(fault), .net(N225), .FEN(FEN[122]), .op(N225_t1) );
fim FAN_N225_2 ( .fault(fault), .net(N225), .FEN(FEN[123]), .op(N225_t2) );
fim FAN_N243_0 ( .fault(fault), .net(N243), .FEN(FEN[124]), .op(N243_t0) );
fim FAN_N243_1 ( .fault(fault), .net(N243), .FEN(FEN[125]), .op(N243_t1) );
fim FAN_N243_2 ( .fault(fault), .net(N243), .FEN(FEN[126]), .op(N243_t2) );
fim FAN_N319_0 ( .fault(fault), .net(N319), .FEN(FEN[127]), .op(N319_t0) );
fim FAN_N319_1 ( .fault(fault), .net(N319), .FEN(FEN[128]), .op(N319_t1) );
fim FAN_N319_2 ( .fault(fault), .net(N319), .FEN(FEN[129]), .op(N319_t2) );
fim FAN_N319_3 ( .fault(fault), .net(N319), .FEN(FEN[130]), .op(N319_t3) );
fim FAN_N319_4 ( .fault(fault), .net(N319), .FEN(FEN[131]), .op(N319_t4) );
fim FAN_N319_5 ( .fault(fault), .net(N319), .FEN(FEN[132]), .op(N319_t5) );
fim FAN_N220_0 ( .fault(fault), .net(N220), .FEN(FEN[133]), .op(N220_t0) );
fim FAN_N220_1 ( .fault(fault), .net(N220), .FEN(FEN[134]), .op(N220_t1) );
fim FAN_N220_2 ( .fault(fault), .net(N220), .FEN(FEN[135]), .op(N220_t2) );
fim FAN_N220_3 ( .fault(fault), .net(N220), .FEN(FEN[136]), .op(N220_t3) );
fim FAN_N229_0 ( .fault(fault), .net(N229), .FEN(FEN[137]), .op(N229_t0) );
fim FAN_N229_1 ( .fault(fault), .net(N229), .FEN(FEN[138]), .op(N229_t1) );
fim FAN_N232_0 ( .fault(fault), .net(N232), .FEN(FEN[139]), .op(N232_t0) );
fim FAN_N232_1 ( .fault(fault), .net(N232), .FEN(FEN[140]), .op(N232_t1) );
fim FAN_N239_0 ( .fault(fault), .net(N239), .FEN(FEN[141]), .op(N239_t0) );
fim FAN_N239_1 ( .fault(fault), .net(N239), .FEN(FEN[142]), .op(N239_t1) );
fim FAN_N239_2 ( .fault(fault), .net(N239), .FEN(FEN[143]), .op(N239_t2) );
fim FAN_N49_0 ( .fault(fault), .net(N49), .FEN(FEN[144]), .op(N49_t0) );
fim FAN_N49_1 ( .fault(fault), .net(N49), .FEN(FEN[145]), .op(N49_t1) );
fim FAN_N49_2 ( .fault(fault), .net(N49), .FEN(FEN[146]), .op(N49_t2) );
fim FAN_N253_0 ( .fault(fault), .net(N253), .FEN(FEN[147]), .op(N253_t0) );
fim FAN_N253_1 ( .fault(fault), .net(N253), .FEN(FEN[148]), .op(N253_t1) );
fim FAN_N247_0 ( .fault(fault), .net(N247), .FEN(FEN[149]), .op(N247_t0) );
fim FAN_N247_1 ( .fault(fault), .net(N247), .FEN(FEN[150]), .op(N247_t1) );
fim FAN_N247_2 ( .fault(fault), .net(N247), .FEN(FEN[151]), .op(N247_t2) );
fim FAN_N326_0 ( .fault(fault), .net(N326), .FEN(FEN[152]), .op(N326_t0) );
fim FAN_N326_1 ( .fault(fault), .net(N326), .FEN(FEN[153]), .op(N326_t1) );
fim FAN_N326_2 ( .fault(fault), .net(N326), .FEN(FEN[154]), .op(N326_t2) );
fim FAN_N326_3 ( .fault(fault), .net(N326), .FEN(FEN[155]), .op(N326_t3) );
fim FAN_N277_0 ( .fault(fault), .net(N277), .FEN(FEN[156]), .op(N277_t0) );
fim FAN_N277_1 ( .fault(fault), .net(N277), .FEN(FEN[157]), .op(N277_t1) );
fim FAN_N280_0 ( .fault(fault), .net(N280), .FEN(FEN[158]), .op(N280_t0) );
fim FAN_N280_1 ( .fault(fault), .net(N280), .FEN(FEN[159]), .op(N280_t1) );
fim FAN_N260_0 ( .fault(fault), .net(N260), .FEN(FEN[160]), .op(N260_t0) );
fim FAN_N260_1 ( .fault(fault), .net(N260), .FEN(FEN[161]), .op(N260_t1) );
fim FAN_N300_0 ( .fault(fault), .net(N300), .FEN(FEN[162]), .op(N300_t0) );
fim FAN_N300_1 ( .fault(fault), .net(N300), .FEN(FEN[163]), .op(N300_t1) );
fim FAN_N201_0 ( .fault(fault), .net(N201), .FEN(FEN[164]), .op(N201_t0) );
fim FAN_N201_1 ( .fault(fault), .net(N201), .FEN(FEN[165]), .op(N201_t1) );
fim FAN_N201_2 ( .fault(fault), .net(N201), .FEN(FEN[166]), .op(N201_t2) );
fim FAN_N201_3 ( .fault(fault), .net(N201), .FEN(FEN[167]), .op(N201_t3) );
fim FAN_N216_0 ( .fault(fault), .net(N216), .FEN(FEN[168]), .op(N216_t0) );
fim FAN_N216_1 ( .fault(fault), .net(N216), .FEN(FEN[169]), .op(N216_t1) );
fim FAN_N216_2 ( .fault(fault), .net(N216), .FEN(FEN[170]), .op(N216_t2) );
fim FAN_N197_0 ( .fault(fault), .net(N197), .FEN(FEN[171]), .op(N197_t0) );
fim FAN_N197_1 ( .fault(fault), .net(N197), .FEN(FEN[172]), .op(N197_t1) );
fim FAN_N197_2 ( .fault(fault), .net(N197), .FEN(FEN[173]), .op(N197_t2) );
fim FAN_N56_0 ( .fault(fault), .net(N56), .FEN(FEN[174]), .op(N56_t0) );
fim FAN_N56_1 ( .fault(fault), .net(N56), .FEN(FEN[175]), .op(N56_t1) );
fim FAN_N56_2 ( .fault(fault), .net(N56), .FEN(FEN[176]), .op(N56_t2) );
fim FAN_N257_0 ( .fault(fault), .net(N257), .FEN(FEN[177]), .op(N257_t0) );
fim FAN_N257_1 ( .fault(fault), .net(N257), .FEN(FEN[178]), .op(N257_t1) );
fim FAN_N235_0 ( .fault(fault), .net(N235), .FEN(FEN[179]), .op(N235_t0) );
fim FAN_N235_1 ( .fault(fault), .net(N235), .FEN(FEN[180]), .op(N235_t1) );
fim FAN_N235_2 ( .fault(fault), .net(N235), .FEN(FEN[181]), .op(N235_t2) );
fim FAN_N60_0 ( .fault(fault), .net(N60), .FEN(FEN[182]), .op(N60_t0) );
fim FAN_N60_1 ( .fault(fault), .net(N60), .FEN(FEN[183]), .op(N60_t1) );
fim FAN_N263_0 ( .fault(fault), .net(N263), .FEN(FEN[184]), .op(N263_t0) );
fim FAN_N263_1 ( .fault(fault), .net(N263), .FEN(FEN[185]), .op(N263_t1) );
fim FAN_N266_0 ( .fault(fault), .net(N266), .FEN(FEN[186]), .op(N266_t0) );
fim FAN_N266_1 ( .fault(fault), .net(N266), .FEN(FEN[187]), .op(N266_t1) );
fim FAN_N269_0 ( .fault(fault), .net(N269), .FEN(FEN[188]), .op(N269_t0) );
fim FAN_N269_1 ( .fault(fault), .net(N269), .FEN(FEN[189]), .op(N269_t1) );
fim FAN_N272_0 ( .fault(fault), .net(N272), .FEN(FEN[190]), .op(N272_t0) );
fim FAN_N272_1 ( .fault(fault), .net(N272), .FEN(FEN[191]), .op(N272_t1) );
fim FAN_N316_0 ( .fault(fault), .net(N316), .FEN(FEN[192]), .op(N316_t0) );
fim FAN_N316_1 ( .fault(fault), .net(N316), .FEN(FEN[193]), .op(N316_t1) );
fim FAN_N212_0 ( .fault(fault), .net(N212), .FEN(FEN[194]), .op(N212_t0) );
fim FAN_N212_1 ( .fault(fault), .net(N212), .FEN(FEN[195]), .op(N212_t1) );
fim FAN_N212_2 ( .fault(fault), .net(N212), .FEN(FEN[196]), .op(N212_t2) );
fim FAN_N53_0 ( .fault(fault), .net(N53), .FEN(FEN[197]), .op(N53_t0) );
fim FAN_N53_1 ( .fault(fault), .net(N53), .FEN(FEN[198]), .op(N53_t1) );
fim FAN_N682_0 ( .fault(fault), .net(N682), .FEN(FEN[199]), .op(N682_t0) );
fim FAN_N682_1 ( .fault(fault), .net(N682), .FEN(FEN[200]), .op(N682_t1) );
fim FAN_N685_0 ( .fault(fault), .net(N685), .FEN(FEN[201]), .op(N685_t0) );
fim FAN_N685_1 ( .fault(fault), .net(N685), .FEN(FEN[202]), .op(N685_t1) );
fim FAN_N616_0 ( .fault(fault), .net(N616), .FEN(FEN[203]), .op(N616_t0) );
fim FAN_N616_1 ( .fault(fault), .net(N616), .FEN(FEN[204]), .op(N616_t1) );
fim FAN_N619_0 ( .fault(fault), .net(N619), .FEN(FEN[205]), .op(N619_t0) );
fim FAN_N619_1 ( .fault(fault), .net(N619), .FEN(FEN[206]), .op(N619_t1) );
fim FAN_N622_0 ( .fault(fault), .net(N622), .FEN(FEN[207]), .op(N622_t0) );
fim FAN_N622_1 ( .fault(fault), .net(N622), .FEN(FEN[208]), .op(N622_t1) );
fim FAN_N625_0 ( .fault(fault), .net(N625), .FEN(FEN[209]), .op(N625_t0) );
fim FAN_N625_1 ( .fault(fault), .net(N625), .FEN(FEN[210]), .op(N625_t1) );
fim FAN_N631_0 ( .fault(fault), .net(N631), .FEN(FEN[211]), .op(N631_t0) );
fim FAN_N631_1 ( .fault(fault), .net(N631), .FEN(FEN[212]), .op(N631_t1) );
fim FAN_N643_0 ( .fault(fault), .net(N643), .FEN(FEN[213]), .op(N643_t0) );
fim FAN_N643_1 ( .fault(fault), .net(N643), .FEN(FEN[214]), .op(N643_t1) );
fim FAN_N649_0 ( .fault(fault), .net(N649), .FEN(FEN[215]), .op(N649_t0) );
fim FAN_N649_1 ( .fault(fault), .net(N649), .FEN(FEN[216]), .op(N649_t1) );
fim FAN_N652_0 ( .fault(fault), .net(N652), .FEN(FEN[217]), .op(N652_t0) );
fim FAN_N652_1 ( .fault(fault), .net(N652), .FEN(FEN[218]), .op(N652_t1) );
fim FAN_N655_0 ( .fault(fault), .net(N655), .FEN(FEN[219]), .op(N655_t0) );
fim FAN_N655_1 ( .fault(fault), .net(N655), .FEN(FEN[220]), .op(N655_t1) );
fim FAN_N612_0 ( .fault(fault), .net(N612), .FEN(FEN[221]), .op(N612_t0) );
fim FAN_N612_1 ( .fault(fault), .net(N612), .FEN(FEN[222]), .op(N612_t1) );
fim FAN_N612_2 ( .fault(fault), .net(N612), .FEN(FEN[223]), .op(N612_t2) );
fim FAN_N608_0 ( .fault(fault), .net(N608), .FEN(FEN[224]), .op(N608_t0) );
fim FAN_N608_1 ( .fault(fault), .net(N608), .FEN(FEN[225]), .op(N608_t1) );
fim FAN_N608_2 ( .fault(fault), .net(N608), .FEN(FEN[226]), .op(N608_t2) );
fim FAN_N661_0 ( .fault(fault), .net(N661), .FEN(FEN[227]), .op(N661_t0) );
fim FAN_N661_1 ( .fault(fault), .net(N661), .FEN(FEN[228]), .op(N661_t1) );
fim FAN_N658_0 ( .fault(fault), .net(N658), .FEN(FEN[229]), .op(N658_t0) );
fim FAN_N658_1 ( .fault(fault), .net(N658), .FEN(FEN[230]), .op(N658_t1) );
fim FAN_N667_0 ( .fault(fault), .net(N667), .FEN(FEN[231]), .op(N667_t0) );
fim FAN_N667_1 ( .fault(fault), .net(N667), .FEN(FEN[232]), .op(N667_t1) );
fim FAN_N664_0 ( .fault(fault), .net(N664), .FEN(FEN[233]), .op(N664_t0) );
fim FAN_N664_1 ( .fault(fault), .net(N664), .FEN(FEN[234]), .op(N664_t1) );
fim FAN_N673_0 ( .fault(fault), .net(N673), .FEN(FEN[235]), .op(N673_t0) );
fim FAN_N673_1 ( .fault(fault), .net(N673), .FEN(FEN[236]), .op(N673_t1) );
fim FAN_N670_0 ( .fault(fault), .net(N670), .FEN(FEN[237]), .op(N670_t0) );
fim FAN_N670_1 ( .fault(fault), .net(N670), .FEN(FEN[238]), .op(N670_t1) );
fim FAN_N679_0 ( .fault(fault), .net(N679), .FEN(FEN[239]), .op(N679_t0) );
fim FAN_N679_1 ( .fault(fault), .net(N679), .FEN(FEN[240]), .op(N679_t1) );
fim FAN_N676_0 ( .fault(fault), .net(N676), .FEN(FEN[241]), .op(N676_t0) );
fim FAN_N676_1 ( .fault(fault), .net(N676), .FEN(FEN[242]), .op(N676_t1) );
fim FAN_N297_0 ( .fault(fault), .net(N297), .FEN(FEN[243]), .op(N297_t0) );
fim FAN_N297_1 ( .fault(fault), .net(N297), .FEN(FEN[244]), .op(N297_t1) );
fim FAN_N603_0 ( .fault(fault), .net(N603), .FEN(FEN[245]), .op(N603_t0) );
fim FAN_N603_1 ( .fault(fault), .net(N603), .FEN(FEN[246]), .op(N603_t1) );
fim FAN_N603_2 ( .fault(fault), .net(N603), .FEN(FEN[247]), .op(N603_t2) );
fim FAN_N603_3 ( .fault(fault), .net(N603), .FEN(FEN[248]), .op(N603_t3) );
fim FAN_N303_0 ( .fault(fault), .net(N303), .FEN(FEN[249]), .op(N303_t0) );
fim FAN_N303_1 ( .fault(fault), .net(N303), .FEN(FEN[250]), .op(N303_t1) );
fim FAN_N338_0 ( .fault(fault), .net(N338), .FEN(FEN[251]), .op(N338_t0) );
fim FAN_N338_1 ( .fault(fault), .net(N338), .FEN(FEN[252]), .op(N338_t1) );
fim FAN_N338_2 ( .fault(fault), .net(N338), .FEN(FEN[253]), .op(N338_t2) );
fim FAN_N338_3 ( .fault(fault), .net(N338), .FEN(FEN[254]), .op(N338_t3) );
fim FAN_N556_0 ( .fault(fault), .net(N556), .FEN(FEN[255]), .op(N556_t0) );
fim FAN_N556_1 ( .fault(fault), .net(N556), .FEN(FEN[256]), .op(N556_t1) );
fim FAN_N688_0 ( .fault(fault), .net(N688), .FEN(FEN[257]), .op(N688_t0) );
fim FAN_N688_1 ( .fault(fault), .net(N688), .FEN(FEN[258]), .op(N688_t1) );
fim FAN_N691_0 ( .fault(fault), .net(N691), .FEN(FEN[259]), .op(N691_t0) );
fim FAN_N691_1 ( .fault(fault), .net(N691), .FEN(FEN[260]), .op(N691_t1) );
fim FAN_N562_0 ( .fault(fault), .net(N562), .FEN(FEN[261]), .op(N562_t0) );
fim FAN_N562_1 ( .fault(fault), .net(N562), .FEN(FEN[262]), .op(N562_t1) );
fim FAN_N694_0 ( .fault(fault), .net(N694), .FEN(FEN[263]), .op(N694_t0) );
fim FAN_N694_1 ( .fault(fault), .net(N694), .FEN(FEN[264]), .op(N694_t1) );
fim FAN_N697_0 ( .fault(fault), .net(N697), .FEN(FEN[265]), .op(N697_t0) );
fim FAN_N697_1 ( .fault(fault), .net(N697), .FEN(FEN[266]), .op(N697_t1) );
fim FAN_N568_0 ( .fault(fault), .net(N568), .FEN(FEN[267]), .op(N568_t0) );
fim FAN_N568_1 ( .fault(fault), .net(N568), .FEN(FEN[268]), .op(N568_t1) );
fim FAN_N700_0 ( .fault(fault), .net(N700), .FEN(FEN[269]), .op(N700_t0) );
fim FAN_N700_1 ( .fault(fault), .net(N700), .FEN(FEN[270]), .op(N700_t1) );
fim FAN_N703_0 ( .fault(fault), .net(N703), .FEN(FEN[271]), .op(N703_t0) );
fim FAN_N703_1 ( .fault(fault), .net(N703), .FEN(FEN[272]), .op(N703_t1) );
fim FAN_N574_0 ( .fault(fault), .net(N574), .FEN(FEN[273]), .op(N574_t0) );
fim FAN_N574_1 ( .fault(fault), .net(N574), .FEN(FEN[274]), .op(N574_t1) );
fim FAN_N580_0 ( .fault(fault), .net(N580), .FEN(FEN[275]), .op(N580_t0) );
fim FAN_N580_1 ( .fault(fault), .net(N580), .FEN(FEN[276]), .op(N580_t1) );
fim FAN_N706_0 ( .fault(fault), .net(N706), .FEN(FEN[277]), .op(N706_t0) );
fim FAN_N706_1 ( .fault(fault), .net(N706), .FEN(FEN[278]), .op(N706_t1) );
fim FAN_N709_0 ( .fault(fault), .net(N709), .FEN(FEN[279]), .op(N709_t0) );
fim FAN_N709_1 ( .fault(fault), .net(N709), .FEN(FEN[280]), .op(N709_t1) );
fim FAN_N586_0 ( .fault(fault), .net(N586), .FEN(FEN[281]), .op(N586_t0) );
fim FAN_N586_1 ( .fault(fault), .net(N586), .FEN(FEN[282]), .op(N586_t1) );
fim FAN_N712_0 ( .fault(fault), .net(N712), .FEN(FEN[283]), .op(N712_t0) );
fim FAN_N712_1 ( .fault(fault), .net(N712), .FEN(FEN[284]), .op(N712_t1) );
fim FAN_N715_0 ( .fault(fault), .net(N715), .FEN(FEN[285]), .op(N715_t0) );
fim FAN_N715_1 ( .fault(fault), .net(N715), .FEN(FEN[286]), .op(N715_t1) );
fim FAN_N592_0 ( .fault(fault), .net(N592), .FEN(FEN[287]), .op(N592_t0) );
fim FAN_N592_1 ( .fault(fault), .net(N592), .FEN(FEN[288]), .op(N592_t1) );
fim FAN_N628_0 ( .fault(fault), .net(N628), .FEN(FEN[289]), .op(N628_t0) );
fim FAN_N628_1 ( .fault(fault), .net(N628), .FEN(FEN[290]), .op(N628_t1) );
fim FAN_N718_0 ( .fault(fault), .net(N718), .FEN(FEN[291]), .op(N718_t0) );
fim FAN_N718_1 ( .fault(fault), .net(N718), .FEN(FEN[292]), .op(N718_t1) );
fim FAN_N721_0 ( .fault(fault), .net(N721), .FEN(FEN[293]), .op(N721_t0) );
fim FAN_N721_1 ( .fault(fault), .net(N721), .FEN(FEN[294]), .op(N721_t1) );
fim FAN_N634_0 ( .fault(fault), .net(N634), .FEN(FEN[295]), .op(N634_t0) );
fim FAN_N634_1 ( .fault(fault), .net(N634), .FEN(FEN[296]), .op(N634_t1) );
fim FAN_N724_0 ( .fault(fault), .net(N724), .FEN(FEN[297]), .op(N724_t0) );
fim FAN_N724_1 ( .fault(fault), .net(N724), .FEN(FEN[298]), .op(N724_t1) );
fim FAN_N727_0 ( .fault(fault), .net(N727), .FEN(FEN[299]), .op(N727_t0) );
fim FAN_N727_1 ( .fault(fault), .net(N727), .FEN(FEN[300]), .op(N727_t1) );
fim FAN_N637_0 ( .fault(fault), .net(N637), .FEN(FEN[301]), .op(N637_t0) );
fim FAN_N637_1 ( .fault(fault), .net(N637), .FEN(FEN[302]), .op(N637_t1) );
fim FAN_N595_0 ( .fault(fault), .net(N595), .FEN(FEN[303]), .op(N595_t0) );
fim FAN_N595_1 ( .fault(fault), .net(N595), .FEN(FEN[304]), .op(N595_t1) );
fim FAN_N730_0 ( .fault(fault), .net(N730), .FEN(FEN[305]), .op(N730_t0) );
fim FAN_N730_1 ( .fault(fault), .net(N730), .FEN(FEN[306]), .op(N730_t1) );
fim FAN_N733_0 ( .fault(fault), .net(N733), .FEN(FEN[307]), .op(N733_t0) );
fim FAN_N733_1 ( .fault(fault), .net(N733), .FEN(FEN[308]), .op(N733_t1) );
fim FAN_N736_0 ( .fault(fault), .net(N736), .FEN(FEN[309]), .op(N736_t0) );
fim FAN_N736_1 ( .fault(fault), .net(N736), .FEN(FEN[310]), .op(N736_t1) );
fim FAN_N739_0 ( .fault(fault), .net(N739), .FEN(FEN[311]), .op(N739_t0) );
fim FAN_N739_1 ( .fault(fault), .net(N739), .FEN(FEN[312]), .op(N739_t1) );
fim FAN_N640_0 ( .fault(fault), .net(N640), .FEN(FEN[313]), .op(N640_t0) );
fim FAN_N640_1 ( .fault(fault), .net(N640), .FEN(FEN[314]), .op(N640_t1) );
fim FAN_N742_0 ( .fault(fault), .net(N742), .FEN(FEN[315]), .op(N742_t0) );
fim FAN_N742_1 ( .fault(fault), .net(N742), .FEN(FEN[316]), .op(N742_t1) );
fim FAN_N745_0 ( .fault(fault), .net(N745), .FEN(FEN[317]), .op(N745_t0) );
fim FAN_N745_1 ( .fault(fault), .net(N745), .FEN(FEN[318]), .op(N745_t1) );
fim FAN_N646_0 ( .fault(fault), .net(N646), .FEN(FEN[319]), .op(N646_t0) );
fim FAN_N646_1 ( .fault(fault), .net(N646), .FEN(FEN[320]), .op(N646_t1) );
fim FAN_N748_0 ( .fault(fault), .net(N748), .FEN(FEN[321]), .op(N748_t0) );
fim FAN_N748_1 ( .fault(fault), .net(N748), .FEN(FEN[322]), .op(N748_t1) );
fim FAN_N751_0 ( .fault(fault), .net(N751), .FEN(FEN[323]), .op(N751_t0) );
fim FAN_N751_1 ( .fault(fault), .net(N751), .FEN(FEN[324]), .op(N751_t1) );
fim FAN_N559_0 ( .fault(fault), .net(N559), .FEN(FEN[325]), .op(N559_t0) );
fim FAN_N559_1 ( .fault(fault), .net(N559), .FEN(FEN[326]), .op(N559_t1) );
fim FAN_N565_0 ( .fault(fault), .net(N565), .FEN(FEN[327]), .op(N565_t0) );
fim FAN_N565_1 ( .fault(fault), .net(N565), .FEN(FEN[328]), .op(N565_t1) );
fim FAN_N571_0 ( .fault(fault), .net(N571), .FEN(FEN[329]), .op(N571_t0) );
fim FAN_N571_1 ( .fault(fault), .net(N571), .FEN(FEN[330]), .op(N571_t1) );
fim FAN_N577_0 ( .fault(fault), .net(N577), .FEN(FEN[331]), .op(N577_t0) );
fim FAN_N577_1 ( .fault(fault), .net(N577), .FEN(FEN[332]), .op(N577_t1) );
fim FAN_N583_0 ( .fault(fault), .net(N583), .FEN(FEN[333]), .op(N583_t0) );
fim FAN_N583_1 ( .fault(fault), .net(N583), .FEN(FEN[334]), .op(N583_t1) );
fim FAN_N589_0 ( .fault(fault), .net(N589), .FEN(FEN[335]), .op(N589_t0) );
fim FAN_N589_1 ( .fault(fault), .net(N589), .FEN(FEN[336]), .op(N589_t1) );
fim FAN_N598_0 ( .fault(fault), .net(N598), .FEN(FEN[337]), .op(N598_t0) );
fim FAN_N598_1 ( .fault(fault), .net(N598), .FEN(FEN[338]), .op(N598_t1) );
fim FAN_N939_0 ( .fault(fault), .net(N939), .FEN(FEN[339]), .op(N939_t0) );
fim FAN_N939_1 ( .fault(fault), .net(N939), .FEN(FEN[340]), .op(N939_t1) );
fim FAN_N935_0 ( .fault(fault), .net(N935), .FEN(FEN[341]), .op(N935_t0) );
fim FAN_N935_1 ( .fault(fault), .net(N935), .FEN(FEN[342]), .op(N935_t1) );
fim FAN_N943_0 ( .fault(fault), .net(N943), .FEN(FEN[343]), .op(N943_t0) );
fim FAN_N943_1 ( .fault(fault), .net(N943), .FEN(FEN[344]), .op(N943_t1) );
fim FAN_N947_0 ( .fault(fault), .net(N947), .FEN(FEN[345]), .op(N947_t0) );
fim FAN_N947_1 ( .fault(fault), .net(N947), .FEN(FEN[346]), .op(N947_t1) );
fim FAN_N955_0 ( .fault(fault), .net(N955), .FEN(FEN[347]), .op(N955_t0) );
fim FAN_N955_1 ( .fault(fault), .net(N955), .FEN(FEN[348]), .op(N955_t1) );
fim FAN_N951_0 ( .fault(fault), .net(N951), .FEN(FEN[349]), .op(N951_t0) );
fim FAN_N951_1 ( .fault(fault), .net(N951), .FEN(FEN[350]), .op(N951_t1) );
fim FAN_N962_0 ( .fault(fault), .net(N962), .FEN(FEN[351]), .op(N962_t0) );
fim FAN_N962_1 ( .fault(fault), .net(N962), .FEN(FEN[352]), .op(N962_t1) );
fim FAN_N969_0 ( .fault(fault), .net(N969), .FEN(FEN[353]), .op(N969_t0) );
fim FAN_N969_1 ( .fault(fault), .net(N969), .FEN(FEN[354]), .op(N969_t1) );
fim FAN_N977_0 ( .fault(fault), .net(N977), .FEN(FEN[355]), .op(N977_t0) );
fim FAN_N977_1 ( .fault(fault), .net(N977), .FEN(FEN[356]), .op(N977_t1) );
fim FAN_N985_0 ( .fault(fault), .net(N985), .FEN(FEN[357]), .op(N985_t0) );
fim FAN_N985_1 ( .fault(fault), .net(N985), .FEN(FEN[358]), .op(N985_t1) );
fim FAN_N998_0 ( .fault(fault), .net(N998), .FEN(FEN[359]), .op(N998_t0) );
fim FAN_N998_1 ( .fault(fault), .net(N998), .FEN(FEN[360]), .op(N998_t1) );
fim FAN_N899_0 ( .fault(fault), .net(N899), .FEN(FEN[361]), .op(N899_t0) );
fim FAN_N899_1 ( .fault(fault), .net(N899), .FEN(FEN[362]), .op(N899_t1) );
fim FAN_N899_2 ( .fault(fault), .net(N899), .FEN(FEN[363]), .op(N899_t2) );
fim FAN_N903_0 ( .fault(fault), .net(N903), .FEN(FEN[364]), .op(N903_t0) );
fim FAN_N903_1 ( .fault(fault), .net(N903), .FEN(FEN[365]), .op(N903_t1) );
fim FAN_N903_2 ( .fault(fault), .net(N903), .FEN(FEN[366]), .op(N903_t2) );
fim FAN_N923_0 ( .fault(fault), .net(N923), .FEN(FEN[367]), .op(N923_t0) );
fim FAN_N923_1 ( .fault(fault), .net(N923), .FEN(FEN[368]), .op(N923_t1) );
fim FAN_N1010_0 ( .fault(fault), .net(N1010), .FEN(FEN[369]), .op(N1010_t0) );
fim FAN_N1010_1 ( .fault(fault), .net(N1010), .FEN(FEN[370]), .op(N1010_t1) );
fim FAN_N1013_0 ( .fault(fault), .net(N1013), .FEN(FEN[371]), .op(N1013_t0) );
fim FAN_N1013_1 ( .fault(fault), .net(N1013), .FEN(FEN[372]), .op(N1013_t1) );
fim FAN_N1016_0 ( .fault(fault), .net(N1016), .FEN(FEN[373]), .op(N1016_t0) );
fim FAN_N1016_1 ( .fault(fault), .net(N1016), .FEN(FEN[374]), .op(N1016_t1) );
fim FAN_N1019_0 ( .fault(fault), .net(N1019), .FEN(FEN[375]), .op(N1019_t0) );
fim FAN_N1019_1 ( .fault(fault), .net(N1019), .FEN(FEN[376]), .op(N1019_t1) );
fim FAN_N1022_0 ( .fault(fault), .net(N1022), .FEN(FEN[377]), .op(N1022_t0) );
fim FAN_N1022_1 ( .fault(fault), .net(N1022), .FEN(FEN[378]), .op(N1022_t1) );
fim FAN_N1025_0 ( .fault(fault), .net(N1025), .FEN(FEN[379]), .op(N1025_t0) );
fim FAN_N1025_1 ( .fault(fault), .net(N1025), .FEN(FEN[380]), .op(N1025_t1) );
fim FAN_N1028_0 ( .fault(fault), .net(N1028), .FEN(FEN[381]), .op(N1028_t0) );
fim FAN_N1028_1 ( .fault(fault), .net(N1028), .FEN(FEN[382]), .op(N1028_t1) );
fim FAN_N959_0 ( .fault(fault), .net(N959), .FEN(FEN[383]), .op(N959_t0) );
fim FAN_N959_1 ( .fault(fault), .net(N959), .FEN(FEN[384]), .op(N959_t1) );
fim FAN_N1031_0 ( .fault(fault), .net(N1031), .FEN(FEN[385]), .op(N1031_t0) );
fim FAN_N1031_1 ( .fault(fault), .net(N1031), .FEN(FEN[386]), .op(N1031_t1) );
fim FAN_N1034_0 ( .fault(fault), .net(N1034), .FEN(FEN[387]), .op(N1034_t0) );
fim FAN_N1034_1 ( .fault(fault), .net(N1034), .FEN(FEN[388]), .op(N1034_t1) );
fim FAN_N965_0 ( .fault(fault), .net(N965), .FEN(FEN[389]), .op(N965_t0) );
fim FAN_N965_1 ( .fault(fault), .net(N965), .FEN(FEN[390]), .op(N965_t1) );
fim FAN_N1037_0 ( .fault(fault), .net(N1037), .FEN(FEN[391]), .op(N1037_t0) );
fim FAN_N1037_1 ( .fault(fault), .net(N1037), .FEN(FEN[392]), .op(N1037_t1) );
fim FAN_N1040_0 ( .fault(fault), .net(N1040), .FEN(FEN[393]), .op(N1040_t0) );
fim FAN_N1040_1 ( .fault(fault), .net(N1040), .FEN(FEN[394]), .op(N1040_t1) );
fim FAN_N973_0 ( .fault(fault), .net(N973), .FEN(FEN[395]), .op(N973_t0) );
fim FAN_N973_1 ( .fault(fault), .net(N973), .FEN(FEN[396]), .op(N973_t1) );
fim FAN_N1043_0 ( .fault(fault), .net(N1043), .FEN(FEN[397]), .op(N1043_t0) );
fim FAN_N1043_1 ( .fault(fault), .net(N1043), .FEN(FEN[398]), .op(N1043_t1) );
fim FAN_N981_0 ( .fault(fault), .net(N981), .FEN(FEN[399]), .op(N981_t0) );
fim FAN_N981_1 ( .fault(fault), .net(N981), .FEN(FEN[400]), .op(N981_t1) );
fim FAN_N1046_0 ( .fault(fault), .net(N1046), .FEN(FEN[401]), .op(N1046_t0) );
fim FAN_N1046_1 ( .fault(fault), .net(N1046), .FEN(FEN[402]), .op(N1046_t1) );
fim FAN_N994_0 ( .fault(fault), .net(N994), .FEN(FEN[403]), .op(N994_t0) );
fim FAN_N994_1 ( .fault(fault), .net(N994), .FEN(FEN[404]), .op(N994_t1) );
fim FAN_N1049_0 ( .fault(fault), .net(N1049), .FEN(FEN[405]), .op(N1049_t0) );
fim FAN_N1049_1 ( .fault(fault), .net(N1049), .FEN(FEN[406]), .op(N1049_t1) );
fim FAN_N907_0 ( .fault(fault), .net(N907), .FEN(FEN[407]), .op(N907_t0) );
fim FAN_N907_1 ( .fault(fault), .net(N907), .FEN(FEN[408]), .op(N907_t1) );
fim FAN_N910_0 ( .fault(fault), .net(N910), .FEN(FEN[409]), .op(N910_t0) );
fim FAN_N910_1 ( .fault(fault), .net(N910), .FEN(FEN[410]), .op(N910_t1) );
fim FAN_N1249_0 ( .fault(fault), .net(N1249), .FEN(FEN[411]), .op(N1249_t0) );
fim FAN_N1249_1 ( .fault(fault), .net(N1249), .FEN(FEN[412]), .op(N1249_t1) );
fim FAN_N1255_0 ( .fault(fault), .net(N1255), .FEN(FEN[413]), .op(N1255_t0) );
fim FAN_N1255_1 ( .fault(fault), .net(N1255), .FEN(FEN[414]), .op(N1255_t1) );
fim FAN_N1252_0 ( .fault(fault), .net(N1252), .FEN(FEN[415]), .op(N1252_t0) );
fim FAN_N1252_1 ( .fault(fault), .net(N1252), .FEN(FEN[416]), .op(N1252_t1) );
fim FAN_N1261_0 ( .fault(fault), .net(N1261), .FEN(FEN[417]), .op(N1261_t0) );
fim FAN_N1261_1 ( .fault(fault), .net(N1261), .FEN(FEN[418]), .op(N1261_t1) );
fim FAN_N1258_0 ( .fault(fault), .net(N1258), .FEN(FEN[419]), .op(N1258_t0) );
fim FAN_N1258_1 ( .fault(fault), .net(N1258), .FEN(FEN[420]), .op(N1258_t1) );
fim FAN_N1232_0 ( .fault(fault), .net(N1232), .FEN(FEN[421]), .op(N1232_t0) );
fim FAN_N1232_1 ( .fault(fault), .net(N1232), .FEN(FEN[422]), .op(N1232_t1) );
fim FAN_N1235_0 ( .fault(fault), .net(N1235), .FEN(FEN[423]), .op(N1235_t0) );
fim FAN_N1235_1 ( .fault(fault), .net(N1235), .FEN(FEN[424]), .op(N1235_t1) );
fim FAN_N1243_0 ( .fault(fault), .net(N1243), .FEN(FEN[425]), .op(N1243_t0) );
fim FAN_N1243_1 ( .fault(fault), .net(N1243), .FEN(FEN[426]), .op(N1243_t1) );
fim FAN_N1246_0 ( .fault(fault), .net(N1246), .FEN(FEN[427]), .op(N1246_t0) );
fim FAN_N1246_1 ( .fault(fault), .net(N1246), .FEN(FEN[428]), .op(N1246_t1) );
fim FAN_N1319_0 ( .fault(fault), .net(N1319), .FEN(FEN[429]), .op(N1319_t0) );
fim FAN_N1319_1 ( .fault(fault), .net(N1319), .FEN(FEN[430]), .op(N1319_t1) );
fim FAN_N1334_0 ( .fault(fault), .net(N1334), .FEN(FEN[431]), .op(N1334_t0) );
fim FAN_N1334_1 ( .fault(fault), .net(N1334), .FEN(FEN[432]), .op(N1334_t1) );
fim FAN_N1264_0 ( .fault(fault), .net(N1264), .FEN(FEN[433]), .op(N1264_t0) );
fim FAN_N1264_1 ( .fault(fault), .net(N1264), .FEN(FEN[434]), .op(N1264_t1) );
fim FAN_N1355_0 ( .fault(fault), .net(N1355), .FEN(FEN[435]), .op(N1355_t0) );
fim FAN_N1355_1 ( .fault(fault), .net(N1355), .FEN(FEN[436]), .op(N1355_t1) );
fim FAN_N1352_0 ( .fault(fault), .net(N1352), .FEN(FEN[437]), .op(N1352_t0) );
fim FAN_N1352_1 ( .fault(fault), .net(N1352), .FEN(FEN[438]), .op(N1352_t1) );
fim FAN_N1358_0 ( .fault(fault), .net(N1358), .FEN(FEN[439]), .op(N1358_t0) );
fim FAN_N1358_1 ( .fault(fault), .net(N1358), .FEN(FEN[440]), .op(N1358_t1) );
fim FAN_N1361_0 ( .fault(fault), .net(N1361), .FEN(FEN[441]), .op(N1361_t0) );
fim FAN_N1361_1 ( .fault(fault), .net(N1361), .FEN(FEN[442]), .op(N1361_t1) );
fim FAN_N1367_0 ( .fault(fault), .net(N1367), .FEN(FEN[443]), .op(N1367_t0) );
fim FAN_N1367_1 ( .fault(fault), .net(N1367), .FEN(FEN[444]), .op(N1367_t1) );
fim FAN_N1364_0 ( .fault(fault), .net(N1364), .FEN(FEN[445]), .op(N1364_t0) );
fim FAN_N1364_1 ( .fault(fault), .net(N1364), .FEN(FEN[446]), .op(N1364_t1) );
fim FAN_N1373_0 ( .fault(fault), .net(N1373), .FEN(FEN[447]), .op(N1373_t0) );
fim FAN_N1373_1 ( .fault(fault), .net(N1373), .FEN(FEN[448]), .op(N1373_t1) );
fim FAN_N1379_0 ( .fault(fault), .net(N1379), .FEN(FEN[449]), .op(N1379_t0) );
fim FAN_N1379_1 ( .fault(fault), .net(N1379), .FEN(FEN[450]), .op(N1379_t1) );
fim FAN_N1383_0 ( .fault(fault), .net(N1383), .FEN(FEN[451]), .op(N1383_t0) );
fim FAN_N1383_1 ( .fault(fault), .net(N1383), .FEN(FEN[452]), .op(N1383_t1) );
fim FAN_N1393_0 ( .fault(fault), .net(N1393), .FEN(FEN[453]), .op(N1393_t0) );
fim FAN_N1393_1 ( .fault(fault), .net(N1393), .FEN(FEN[454]), .op(N1393_t1) );
fim FAN_N1370_0 ( .fault(fault), .net(N1370), .FEN(FEN[455]), .op(N1370_t0) );
fim FAN_N1370_1 ( .fault(fault), .net(N1370), .FEN(FEN[456]), .op(N1370_t1) );
fim FAN_N1376_0 ( .fault(fault), .net(N1376), .FEN(FEN[457]), .op(N1376_t0) );
fim FAN_N1376_1 ( .fault(fault), .net(N1376), .FEN(FEN[458]), .op(N1376_t1) );
fim FAN_N1390_0 ( .fault(fault), .net(N1390), .FEN(FEN[459]), .op(N1390_t0) );
fim FAN_N1390_1 ( .fault(fault), .net(N1390), .FEN(FEN[460]), .op(N1390_t1) );
fim FAN_N1419_0 ( .fault(fault), .net(N1419), .FEN(FEN[461]), .op(N1419_t0) );
fim FAN_N1419_1 ( .fault(fault), .net(N1419), .FEN(FEN[462]), .op(N1419_t1) );
fim FAN_N1416_0 ( .fault(fault), .net(N1416), .FEN(FEN[463]), .op(N1416_t0) );
fim FAN_N1416_1 ( .fault(fault), .net(N1416), .FEN(FEN[464]), .op(N1416_t1) );
fim FAN_N1440_0 ( .fault(fault), .net(N1440), .FEN(FEN[465]), .op(N1440_t0) );
fim FAN_N1440_1 ( .fault(fault), .net(N1440), .FEN(FEN[466]), .op(N1440_t1) );
fim FAN_N1472_0 ( .fault(fault), .net(N1472), .FEN(FEN[467]), .op(N1472_t0) );
fim FAN_N1472_1 ( .fault(fault), .net(N1472), .FEN(FEN[468]), .op(N1472_t1) );
fim FAN_N1478_0 ( .fault(fault), .net(N1478), .FEN(FEN[469]), .op(N1478_t0) );
fim FAN_N1478_1 ( .fault(fault), .net(N1478), .FEN(FEN[470]), .op(N1478_t1) );
fim FAN_N1481_0 ( .fault(fault), .net(N1481), .FEN(FEN[471]), .op(N1481_t0) );
fim FAN_N1481_1 ( .fault(fault), .net(N1481), .FEN(FEN[472]), .op(N1481_t1) );
fim FAN_N1484_0 ( .fault(fault), .net(N1484), .FEN(FEN[473]), .op(N1484_t0) );
fim FAN_N1484_1 ( .fault(fault), .net(N1484), .FEN(FEN[474]), .op(N1484_t1) );
fim FAN_N1510_0 ( .fault(fault), .net(N1510), .FEN(FEN[475]), .op(N1510_t0) );
fim FAN_N1510_1 ( .fault(fault), .net(N1510), .FEN(FEN[476]), .op(N1510_t1) );
fim FAN_N1522_0 ( .fault(fault), .net(N1522), .FEN(FEN[477]), .op(N1522_t0) );
fim FAN_N1522_1 ( .fault(fault), .net(N1522), .FEN(FEN[478]), .op(N1522_t1) );
fim FAN_N1522_2 ( .fault(fault), .net(N1522), .FEN(FEN[479]), .op(N1522_t2) );
fim FAN_N1534_0 ( .fault(fault), .net(N1534), .FEN(FEN[480]), .op(N1534_t0) );
fim FAN_N1534_1 ( .fault(fault), .net(N1534), .FEN(FEN[481]), .op(N1534_t1) );
fim FAN_N1537_0 ( .fault(fault), .net(N1537), .FEN(FEN[482]), .op(N1537_t0) );
fim FAN_N1537_1 ( .fault(fault), .net(N1537), .FEN(FEN[483]), .op(N1537_t1) );
fim FAN_N1540_0 ( .fault(fault), .net(N1540), .FEN(FEN[484]), .op(N1540_t0) );
fim FAN_N1540_1 ( .fault(fault), .net(N1540), .FEN(FEN[485]), .op(N1540_t1) );
fim FAN_N1517_0 ( .fault(fault), .net(N1517), .FEN(FEN[486]), .op(N1517_t0) );
fim FAN_N1517_1 ( .fault(fault), .net(N1517), .FEN(FEN[487]), .op(N1517_t1) );
fim FAN_N1514_0 ( .fault(fault), .net(N1514), .FEN(FEN[488]), .op(N1514_t0) );
fim FAN_N1514_1 ( .fault(fault), .net(N1514), .FEN(FEN[489]), .op(N1514_t1) );
fim FAN_N1557_0 ( .fault(fault), .net(N1557), .FEN(FEN[490]), .op(N1557_t0) );
fim FAN_N1557_1 ( .fault(fault), .net(N1557), .FEN(FEN[491]), .op(N1557_t1) );
fim FAN_N1557_2 ( .fault(fault), .net(N1557), .FEN(FEN[492]), .op(N1557_t2) );
fim FAN_N1554_0 ( .fault(fault), .net(N1554), .FEN(FEN[493]), .op(N1554_t0) );
fim FAN_N1554_1 ( .fault(fault), .net(N1554), .FEN(FEN[494]), .op(N1554_t1) );
fim FAN_N1571_0 ( .fault(fault), .net(N1571), .FEN(FEN[495]), .op(N1571_t0) );
fim FAN_N1571_1 ( .fault(fault), .net(N1571), .FEN(FEN[496]), .op(N1571_t1) );
fim FAN_N1576_0 ( .fault(fault), .net(N1576), .FEN(FEN[497]), .op(N1576_t0) );
fim FAN_N1576_1 ( .fault(fault), .net(N1576), .FEN(FEN[498]), .op(N1576_t1) );
fim FAN_N1561_0 ( .fault(fault), .net(N1561), .FEN(FEN[499]), .op(N1561_t0) );
fim FAN_N1561_1 ( .fault(fault), .net(N1561), .FEN(FEN[500]), .op(N1561_t1) );
fim FAN_N1546_0 ( .fault(fault), .net(N1546), .FEN(FEN[501]), .op(N1546_t0) );
fim FAN_N1546_1 ( .fault(fault), .net(N1546), .FEN(FEN[502]), .op(N1546_t1) );
fim FAN_N1596_0 ( .fault(fault), .net(N1596), .FEN(FEN[503]), .op(N1596_t0) );
fim FAN_N1596_1 ( .fault(fault), .net(N1596), .FEN(FEN[504]), .op(N1596_t1) );
fim FAN_N1600_0 ( .fault(fault), .net(N1600), .FEN(FEN[505]), .op(N1600_t0) );
fim FAN_N1600_1 ( .fault(fault), .net(N1600), .FEN(FEN[506]), .op(N1600_t1) );
fim FAN_N1603_0 ( .fault(fault), .net(N1603), .FEN(FEN[507]), .op(N1603_t0) );
fim FAN_N1603_1 ( .fault(fault), .net(N1603), .FEN(FEN[508]), .op(N1603_t1) );
fim FAN_N1606_0 ( .fault(fault), .net(N1606), .FEN(FEN[509]), .op(N1606_t0) );
fim FAN_N1606_1 ( .fault(fault), .net(N1606), .FEN(FEN[510]), .op(N1606_t1) );
fim FAN_N1609_0 ( .fault(fault), .net(N1609), .FEN(FEN[511]), .op(N1609_t0) );
fim FAN_N1609_1 ( .fault(fault), .net(N1609), .FEN(FEN[512]), .op(N1609_t1) );
fim FAN_N1612_0 ( .fault(fault), .net(N1612), .FEN(FEN[513]), .op(N1612_t0) );
fim FAN_N1612_1 ( .fault(fault), .net(N1612), .FEN(FEN[514]), .op(N1612_t1) );
fim FAN_N1615_0 ( .fault(fault), .net(N1615), .FEN(FEN[515]), .op(N1615_t0) );
fim FAN_N1615_1 ( .fault(fault), .net(N1615), .FEN(FEN[516]), .op(N1615_t1) );
fim FAN_N1588_0 ( .fault(fault), .net(N1588), .FEN(FEN[517]), .op(N1588_t0) );
fim FAN_N1588_1 ( .fault(fault), .net(N1588), .FEN(FEN[518]), .op(N1588_t1) );
fim FAN_N1643_0 ( .fault(fault), .net(N1643), .FEN(FEN[519]), .op(N1643_t0) );
fim FAN_N1643_1 ( .fault(fault), .net(N1643), .FEN(FEN[520]), .op(N1643_t1) );
fim FAN_N1647_0 ( .fault(fault), .net(N1647), .FEN(FEN[521]), .op(N1647_t0) );
fim FAN_N1647_1 ( .fault(fault), .net(N1647), .FEN(FEN[522]), .op(N1647_t1) );
fim FAN_N1651_0 ( .fault(fault), .net(N1651), .FEN(FEN[523]), .op(N1651_t0) );
fim FAN_N1651_1 ( .fault(fault), .net(N1651), .FEN(FEN[524]), .op(N1651_t1) );
fim FAN_N1620_0 ( .fault(fault), .net(N1620), .FEN(FEN[525]), .op(N1620_t0) );
fim FAN_N1620_1 ( .fault(fault), .net(N1620), .FEN(FEN[526]), .op(N1620_t1) );
fim FAN_N1658_0 ( .fault(fault), .net(N1658), .FEN(FEN[527]), .op(N1658_t0) );
fim FAN_N1658_1 ( .fault(fault), .net(N1658), .FEN(FEN[528]), .op(N1658_t1) );
fim FAN_N1661_0 ( .fault(fault), .net(N1661), .FEN(FEN[529]), .op(N1661_t0) );
fim FAN_N1661_1 ( .fault(fault), .net(N1661), .FEN(FEN[530]), .op(N1661_t1) );
fim FAN_N1640_0 ( .fault(fault), .net(N1640), .FEN(FEN[531]), .op(N1640_t0) );
fim FAN_N1640_1 ( .fault(fault), .net(N1640), .FEN(FEN[532]), .op(N1640_t1) );
fim FAN_N1664_0 ( .fault(fault), .net(N1664), .FEN(FEN[533]), .op(N1664_t0) );
fim FAN_N1664_1 ( .fault(fault), .net(N1664), .FEN(FEN[534]), .op(N1664_t1) );
fim FAN_N1623_0 ( .fault(fault), .net(N1623), .FEN(FEN[535]), .op(N1623_t0) );
fim FAN_N1623_1 ( .fault(fault), .net(N1623), .FEN(FEN[536]), .op(N1623_t1) );
fim FAN_N1685_0 ( .fault(fault), .net(N1685), .FEN(FEN[537]), .op(N1685_t0) );
fim FAN_N1685_1 ( .fault(fault), .net(N1685), .FEN(FEN[538]), .op(N1685_t1) );
fim FAN_N1697_0 ( .fault(fault), .net(N1697), .FEN(FEN[539]), .op(N1697_t0) );
fim FAN_N1697_1 ( .fault(fault), .net(N1697), .FEN(FEN[540]), .op(N1697_t1) );
fim FAN_N1701_0 ( .fault(fault), .net(N1701), .FEN(FEN[541]), .op(N1701_t0) );
fim FAN_N1701_1 ( .fault(fault), .net(N1701), .FEN(FEN[542]), .op(N1701_t1) );
fim FAN_N1717_0 ( .fault(fault), .net(N1717), .FEN(FEN[543]), .op(N1717_t0) );
fim FAN_N1717_1 ( .fault(fault), .net(N1717), .FEN(FEN[544]), .op(N1717_t1) );
fim FAN_N1723_0 ( .fault(fault), .net(N1723), .FEN(FEN[545]), .op(N1723_t0) );
fim FAN_N1723_1 ( .fault(fault), .net(N1723), .FEN(FEN[546]), .op(N1723_t1) );
fim FAN_N1731_0 ( .fault(fault), .net(N1731), .FEN(FEN[547]), .op(N1731_t0) );
fim FAN_N1731_1 ( .fault(fault), .net(N1731), .FEN(FEN[548]), .op(N1731_t1) );
fim FAN_N1714_0 ( .fault(fault), .net(N1714), .FEN(FEN[549]), .op(N1714_t0) );
fim FAN_N1714_1 ( .fault(fault), .net(N1714), .FEN(FEN[550]), .op(N1714_t1) );
fim FAN_N1734_0 ( .fault(fault), .net(N1734), .FEN(FEN[551]), .op(N1734_t0) );
fim FAN_N1734_1 ( .fault(fault), .net(N1734), .FEN(FEN[552]), .op(N1734_t1) );
fim FAN_N1751_0 ( .fault(fault), .net(N1751), .FEN(FEN[553]), .op(N1751_t0) );
fim FAN_N1751_1 ( .fault(fault), .net(N1751), .FEN(FEN[554]), .op(N1751_t1) );
fim FAN_N1742_0 ( .fault(fault), .net(N1742), .FEN(FEN[555]), .op(N1742_t0) );
fim FAN_N1742_1 ( .fault(fault), .net(N1742), .FEN(FEN[556]), .op(N1742_t1) );
fim FAN_N290_0 ( .fault(fault), .net(N290), .FEN(FEN[557]), .op(N290_t0) );
fim FAN_N290_1 ( .fault(fault), .net(N290), .FEN(FEN[558]), .op(N290_t1) );
fim FAN_N290_2 ( .fault(fault), .net(N290), .FEN(FEN[559]), .op(N290_t2) );
fim FAN_N290_3 ( .fault(fault), .net(N290), .FEN(FEN[560]), .op(N290_t3) );
fim FAN_N290_4 ( .fault(fault), .net(N290), .FEN(FEN[561]), .op(N290_t4) );
fim FAN_N290_5 ( .fault(fault), .net(N290), .FEN(FEN[562]), .op(N290_t5) );
fim FAN_N1748_0 ( .fault(fault), .net(N1748), .FEN(FEN[563]), .op(N1748_t0) );
fim FAN_N1748_1 ( .fault(fault), .net(N1748), .FEN(FEN[564]), .op(N1748_t1) );
fim FAN_N1777_0 ( .fault(fault), .net(N1777), .FEN(FEN[565]), .op(N1777_t0) );
fim FAN_N1777_1 ( .fault(fault), .net(N1777), .FEN(FEN[566]), .op(N1777_t1) );
fim FAN_N1774_0 ( .fault(fault), .net(N1774), .FEN(FEN[567]), .op(N1774_t0) );
fim FAN_N1774_1 ( .fault(fault), .net(N1774), .FEN(FEN[568]), .op(N1774_t1) );
fim FAN_N1788_0 ( .fault(fault), .net(N1788), .FEN(FEN[569]), .op(N1788_t0) );
fim FAN_N1788_1 ( .fault(fault), .net(N1788), .FEN(FEN[570]), .op(N1788_t1) );
fim FAN_N1815_0 ( .fault(fault), .net(N1815), .FEN(FEN[571]), .op(N1815_t0) );
fim FAN_N1815_1 ( .fault(fault), .net(N1815), .FEN(FEN[572]), .op(N1815_t1) );
fim FAN_N1818_0 ( .fault(fault), .net(N1818), .FEN(FEN[573]), .op(N1818_t0) );
fim FAN_N1818_1 ( .fault(fault), .net(N1818), .FEN(FEN[574]), .op(N1818_t1) );
fim FAN_N1798_0 ( .fault(fault), .net(N1798), .FEN(FEN[575]), .op(N1798_t0) );
fim FAN_N1798_1 ( .fault(fault), .net(N1798), .FEN(FEN[576]), .op(N1798_t1) );
fim FAN_N1812_0 ( .fault(fault), .net(N1812), .FEN(FEN[577]), .op(N1812_t0) );
fim FAN_N1812_1 ( .fault(fault), .net(N1812), .FEN(FEN[578]), .op(N1812_t1) );
fim FAN_N1802_0 ( .fault(fault), .net(N1802), .FEN(FEN[579]), .op(N1802_t0) );
fim FAN_N1802_1 ( .fault(fault), .net(N1802), .FEN(FEN[580]), .op(N1802_t1) );
fim FAN_N1841_0 ( .fault(fault), .net(N1841), .FEN(FEN[581]), .op(N1841_t0) );
fim FAN_N1841_1 ( .fault(fault), .net(N1841), .FEN(FEN[582]), .op(N1841_t1) );
fim FAN_N1830_0 ( .fault(fault), .net(N1830), .FEN(FEN[583]), .op(N1830_t0) );
fim FAN_N1830_1 ( .fault(fault), .net(N1830), .FEN(FEN[584]), .op(N1830_t1) );
fim FAN_N1838_0 ( .fault(fault), .net(N1838), .FEN(FEN[585]), .op(N1838_t0) );
fim FAN_N1838_1 ( .fault(fault), .net(N1838), .FEN(FEN[586]), .op(N1838_t1) );
fim FAN_N1866_0 ( .fault(fault), .net(N1866), .FEN(FEN[587]), .op(N1866_t0) );
fim FAN_N1866_1 ( .fault(fault), .net(N1866), .FEN(FEN[588]), .op(N1866_t1) );
fim FAN_N1872_0 ( .fault(fault), .net(N1872), .FEN(FEN[589]), .op(N1872_t0) );
fim FAN_N1872_1 ( .fault(fault), .net(N1872), .FEN(FEN[590]), .op(N1872_t1) );
fim FAN_N1869_0 ( .fault(fault), .net(N1869), .FEN(FEN[591]), .op(N1869_t0) );
fim FAN_N1869_1 ( .fault(fault), .net(N1869), .FEN(FEN[592]), .op(N1869_t1) );
fim FAN_N1875_0 ( .fault(fault), .net(N1875), .FEN(FEN[593]), .op(N1875_t0) );
fim FAN_N1875_1 ( .fault(fault), .net(N1875), .FEN(FEN[594]), .op(N1875_t1) );
fim FAN_N1858_0 ( .fault(fault), .net(N1858), .FEN(FEN[595]), .op(N1858_t0) );
fim FAN_N1858_1 ( .fault(fault), .net(N1858), .FEN(FEN[596]), .op(N1858_t1) );
fim FAN_N1898_0 ( .fault(fault), .net(N1898), .FEN(FEN[597]), .op(N1898_t0) );
fim FAN_N1898_1 ( .fault(fault), .net(N1898), .FEN(FEN[598]), .op(N1898_t1) );
fim FAN_N1902_0 ( .fault(fault), .net(N1902), .FEN(FEN[599]), .op(N1902_t0) );
fim FAN_N1902_1 ( .fault(fault), .net(N1902), .FEN(FEN[600]), .op(N1902_t1) );
fim FAN_N1879_0 ( .fault(fault), .net(N1879), .FEN(FEN[601]), .op(N1879_t0) );
fim FAN_N1879_1 ( .fault(fault), .net(N1879), .FEN(FEN[602]), .op(N1879_t1) );
fim FAN_N1889_0 ( .fault(fault), .net(N1889), .FEN(FEN[603]), .op(N1889_t0) );
fim FAN_N1889_1 ( .fault(fault), .net(N1889), .FEN(FEN[604]), .op(N1889_t1) );
fim FAN_N1930_0 ( .fault(fault), .net(N1930), .FEN(FEN[605]), .op(N1930_t0) );
fim FAN_N1930_1 ( .fault(fault), .net(N1930), .FEN(FEN[606]), .op(N1930_t1) );
fim FAN_N1927_0 ( .fault(fault), .net(N1927), .FEN(FEN[607]), .op(N1927_t0) );
fim FAN_N1927_1 ( .fault(fault), .net(N1927), .FEN(FEN[608]), .op(N1927_t1) );
fim FAN_N1933_0 ( .fault(fault), .net(N1933), .FEN(FEN[609]), .op(N1933_t0) );
fim FAN_N1933_1 ( .fault(fault), .net(N1933), .FEN(FEN[610]), .op(N1933_t1) );
fim FAN_N1944_0 ( .fault(fault), .net(N1944), .FEN(FEN[611]), .op(N1944_t0) );
fim FAN_N1944_1 ( .fault(fault), .net(N1944), .FEN(FEN[612]), .op(N1944_t1) );
fim FAN_N1947_0 ( .fault(fault), .net(N1947), .FEN(FEN[613]), .op(N1947_t0) );
fim FAN_N1947_1 ( .fault(fault), .net(N1947), .FEN(FEN[614]), .op(N1947_t1) );
fim FAN_N1953_0 ( .fault(fault), .net(N1953), .FEN(FEN[615]), .op(N1953_t0) );
fim FAN_N1953_1 ( .fault(fault), .net(N1953), .FEN(FEN[616]), .op(N1953_t1) );
fim FAN_N1950_0 ( .fault(fault), .net(N1950), .FEN(FEN[617]), .op(N1950_t0) );
fim FAN_N1950_1 ( .fault(fault), .net(N1950), .FEN(FEN[618]), .op(N1950_t1) );
fim FAN_N1958_0 ( .fault(fault), .net(N1958), .FEN(FEN[619]), .op(N1958_t0) );
fim FAN_N1958_1 ( .fault(fault), .net(N1958), .FEN(FEN[620]), .op(N1958_t1) );
fim FAN_N1961_0 ( .fault(fault), .net(N1961), .FEN(FEN[621]), .op(N1961_t0) );
fim FAN_N1961_1 ( .fault(fault), .net(N1961), .FEN(FEN[622]), .op(N1961_t1) );
fim FAN_N1965_0 ( .fault(fault), .net(N1965), .FEN(FEN[623]), .op(N1965_t0) );
fim FAN_N1965_1 ( .fault(fault), .net(N1965), .FEN(FEN[624]), .op(N1965_t1) );
fim FAN_N1968_0 ( .fault(fault), .net(N1968), .FEN(FEN[625]), .op(N1968_t0) );
fim FAN_N1968_1 ( .fault(fault), .net(N1968), .FEN(FEN[626]), .op(N1968_t1) );
fim FAN_N1987_0 ( .fault(fault), .net(N1987), .FEN(FEN[627]), .op(N1987_t0) );
fim FAN_N1987_1 ( .fault(fault), .net(N1987), .FEN(FEN[628]), .op(N1987_t1) );
fim FAN_N1980_0 ( .fault(fault), .net(N1980), .FEN(FEN[629]), .op(N1980_t0) );
fim FAN_N1980_1 ( .fault(fault), .net(N1980), .FEN(FEN[630]), .op(N1980_t1) );
fim FAN_N2027_0 ( .fault(fault), .net(N2027), .FEN(FEN[631]), .op(N2027_t0) );
fim FAN_N2027_1 ( .fault(fault), .net(N2027), .FEN(FEN[632]), .op(N2027_t1) );
fim FAN_N2052_0 ( .fault(fault), .net(N2052), .FEN(FEN[633]), .op(N2052_t0) );
fim FAN_N2052_1 ( .fault(fault), .net(N2052), .FEN(FEN[634]), .op(N2052_t1) );
fim FAN_N2055_0 ( .fault(fault), .net(N2055), .FEN(FEN[635]), .op(N2055_t0) );
fim FAN_N2055_1 ( .fault(fault), .net(N2055), .FEN(FEN[636]), .op(N2055_t1) );
fim FAN_N2042_0 ( .fault(fault), .net(N2042), .FEN(FEN[637]), .op(N2042_t0) );
fim FAN_N2042_1 ( .fault(fault), .net(N2042), .FEN(FEN[638]), .op(N2042_t1) );
fim FAN_N2030_0 ( .fault(fault), .net(N2030), .FEN(FEN[639]), .op(N2030_t0) );
fim FAN_N2030_1 ( .fault(fault), .net(N2030), .FEN(FEN[640]), .op(N2030_t1) );
fim FAN_N2068_0 ( .fault(fault), .net(N2068), .FEN(FEN[641]), .op(N2068_t0) );
fim FAN_N2068_1 ( .fault(fault), .net(N2068), .FEN(FEN[642]), .op(N2068_t1) );
fim FAN_N2033_0 ( .fault(fault), .net(N2033), .FEN(FEN[643]), .op(N2033_t0) );
fim FAN_N2033_1 ( .fault(fault), .net(N2033), .FEN(FEN[644]), .op(N2033_t1) );
fim FAN_N2071_0 ( .fault(fault), .net(N2071), .FEN(FEN[645]), .op(N2071_t0) );
fim FAN_N2071_1 ( .fault(fault), .net(N2071), .FEN(FEN[646]), .op(N2071_t1) );
fim FAN_N2062_0 ( .fault(fault), .net(N2062), .FEN(FEN[647]), .op(N2062_t0) );
fim FAN_N2062_1 ( .fault(fault), .net(N2062), .FEN(FEN[648]), .op(N2062_t1) );
fim FAN_N2078_0 ( .fault(fault), .net(N2078), .FEN(FEN[649]), .op(N2078_t0) );
fim FAN_N2078_1 ( .fault(fault), .net(N2078), .FEN(FEN[650]), .op(N2078_t1) );
fim FAN_N2081_0 ( .fault(fault), .net(N2081), .FEN(FEN[651]), .op(N2081_t0) );
fim FAN_N2081_1 ( .fault(fault), .net(N2081), .FEN(FEN[652]), .op(N2081_t1) );
fim FAN_N2151_0 ( .fault(fault), .net(N2151), .FEN(FEN[653]), .op(N2151_t0) );
fim FAN_N2151_1 ( .fault(fault), .net(N2151), .FEN(FEN[654]), .op(N2151_t1) );
fim FAN_N2148_0 ( .fault(fault), .net(N2148), .FEN(FEN[655]), .op(N2148_t0) );
fim FAN_N2148_1 ( .fault(fault), .net(N2148), .FEN(FEN[656]), .op(N2148_t1) );
fim FAN_N2199_0 ( .fault(fault), .net(N2199), .FEN(FEN[657]), .op(N2199_t0) );
fim FAN_N2199_1 ( .fault(fault), .net(N2199), .FEN(FEN[658]), .op(N2199_t1) );
fim FAN_N2196_0 ( .fault(fault), .net(N2196), .FEN(FEN[659]), .op(N2196_t0) );
fim FAN_N2196_1 ( .fault(fault), .net(N2196), .FEN(FEN[660]), .op(N2196_t1) );
fim FAN_N2205_0 ( .fault(fault), .net(N2205), .FEN(FEN[661]), .op(N2205_t0) );
fim FAN_N2205_1 ( .fault(fault), .net(N2205), .FEN(FEN[662]), .op(N2205_t1) );
fim FAN_N2202_0 ( .fault(fault), .net(N2202), .FEN(FEN[663]), .op(N2202_t0) );
fim FAN_N2202_1 ( .fault(fault), .net(N2202), .FEN(FEN[664]), .op(N2202_t1) );
fim FAN_N2237_0 ( .fault(fault), .net(N2237), .FEN(FEN[665]), .op(N2237_t0) );
fim FAN_N2237_1 ( .fault(fault), .net(N2237), .FEN(FEN[666]), .op(N2237_t1) );
fim FAN_N2241_0 ( .fault(fault), .net(N2241), .FEN(FEN[667]), .op(N2241_t0) );
fim FAN_N2241_1 ( .fault(fault), .net(N2241), .FEN(FEN[668]), .op(N2241_t1) );
fim FAN_N1164_0 ( .fault(fault), .net(N1164), .FEN(FEN[669]), .op(N1164_t0) );
fim FAN_N1164_1 ( .fault(fault), .net(N1164), .FEN(FEN[670]), .op(N1164_t1) );
fim FAN_N2245_0 ( .fault(fault), .net(N2245), .FEN(FEN[671]), .op(N2245_t0) );
fim FAN_N2245_1 ( .fault(fault), .net(N2245), .FEN(FEN[672]), .op(N2245_t1) );
fim FAN_N1168_0 ( .fault(fault), .net(N1168), .FEN(FEN[673]), .op(N1168_t0) );
fim FAN_N1168_1 ( .fault(fault), .net(N1168), .FEN(FEN[674]), .op(N1168_t1) );
fim FAN_N2266_0 ( .fault(fault), .net(N2266), .FEN(FEN[675]), .op(N2266_t0) );
fim FAN_N2266_1 ( .fault(fault), .net(N2266), .FEN(FEN[676]), .op(N2266_t1) );
fim FAN_N2272_0 ( .fault(fault), .net(N2272), .FEN(FEN[677]), .op(N2272_t0) );
fim FAN_N2272_1 ( .fault(fault), .net(N2272), .FEN(FEN[678]), .op(N2272_t1) );
fim FAN_N2086_0 ( .fault(fault), .net(N2086), .FEN(FEN[679]), .op(N2086_t0) );
fim FAN_N2086_1 ( .fault(fault), .net(N2086), .FEN(FEN[680]), .op(N2086_t1) );
fim FAN_N2257_0 ( .fault(fault), .net(N2257), .FEN(FEN[681]), .op(N2257_t0) );
fim FAN_N2257_1 ( .fault(fault), .net(N2257), .FEN(FEN[682]), .op(N2257_t1) );
fim FAN_N2089_0 ( .fault(fault), .net(N2089), .FEN(FEN[683]), .op(N2089_t0) );
fim FAN_N2089_1 ( .fault(fault), .net(N2089), .FEN(FEN[684]), .op(N2089_t1) );
fim FAN_N2260_0 ( .fault(fault), .net(N2260), .FEN(FEN[685]), .op(N2260_t0) );
fim FAN_N2260_1 ( .fault(fault), .net(N2260), .FEN(FEN[686]), .op(N2260_t1) );
fim FAN_N2279_0 ( .fault(fault), .net(N2279), .FEN(FEN[687]), .op(N2279_t0) );
fim FAN_N2279_1 ( .fault(fault), .net(N2279), .FEN(FEN[688]), .op(N2279_t1) );
fim FAN_N313_0 ( .fault(fault), .net(N313), .FEN(FEN[689]), .op(N313_t0) );
fim FAN_N313_1 ( .fault(fault), .net(N313), .FEN(FEN[690]), .op(N313_t1) );
fim FAN_N2263_0 ( .fault(fault), .net(N2263), .FEN(FEN[691]), .op(N2263_t0) );
fim FAN_N2263_1 ( .fault(fault), .net(N2263), .FEN(FEN[692]), .op(N2263_t1) );
fim FAN_N2269_0 ( .fault(fault), .net(N2269), .FEN(FEN[693]), .op(N2269_t0) );
fim FAN_N2269_1 ( .fault(fault), .net(N2269), .FEN(FEN[694]), .op(N2269_t1) );
fim FAN_N2286_0 ( .fault(fault), .net(N2286), .FEN(FEN[695]), .op(N2286_t0) );
fim FAN_N2286_1 ( .fault(fault), .net(N2286), .FEN(FEN[696]), .op(N2286_t1) );
fim FAN_N2286_2 ( .fault(fault), .net(N2286), .FEN(FEN[697]), .op(N2286_t2) );
fim FAN_N2286_3 ( .fault(fault), .net(N2286), .FEN(FEN[698]), .op(N2286_t3) );
fim FAN_N2286_4 ( .fault(fault), .net(N2286), .FEN(FEN[699]), .op(N2286_t4) );
fim FAN_N2286_5 ( .fault(fault), .net(N2286), .FEN(FEN[700]), .op(N2286_t5) );
fim FAN_N2286_6 ( .fault(fault), .net(N2286), .FEN(FEN[701]), .op(N2286_t6) );
fim FAN_N2286_7 ( .fault(fault), .net(N2286), .FEN(FEN[702]), .op(N2286_t7) );
fim FAN_N2286_8 ( .fault(fault), .net(N2286), .FEN(FEN[703]), .op(N2286_t8) );
fim FAN_N2286_9 ( .fault(fault), .net(N2286), .FEN(FEN[704]), .op(N2286_t9) );
fim FAN_N2315_0 ( .fault(fault), .net(N2315), .FEN(FEN[705]), .op(N2315_t0) );
fim FAN_N2315_1 ( .fault(fault), .net(N2315), .FEN(FEN[706]), .op(N2315_t1) );
fim FAN_N2315_2 ( .fault(fault), .net(N2315), .FEN(FEN[707]), .op(N2315_t2) );
fim FAN_N2315_3 ( .fault(fault), .net(N2315), .FEN(FEN[708]), .op(N2315_t3) );
fim FAN_N2315_4 ( .fault(fault), .net(N2315), .FEN(FEN[709]), .op(N2315_t4) );
fim FAN_N2315_5 ( .fault(fault), .net(N2315), .FEN(FEN[710]), .op(N2315_t5) );
fim FAN_N2315_6 ( .fault(fault), .net(N2315), .FEN(FEN[711]), .op(N2315_t6) );
fim FAN_N2315_7 ( .fault(fault), .net(N2315), .FEN(FEN[712]), .op(N2315_t7) );
fim FAN_N2315_8 ( .fault(fault), .net(N2315), .FEN(FEN[713]), .op(N2315_t8) );
fim FAN_N2315_9 ( .fault(fault), .net(N2315), .FEN(FEN[714]), .op(N2315_t9) );
fim FAN_N2361_0 ( .fault(fault), .net(N2361), .FEN(FEN[715]), .op(N2361_t0) );
fim FAN_N2361_1 ( .fault(fault), .net(N2361), .FEN(FEN[716]), .op(N2361_t1) );
fim FAN_N2361_2 ( .fault(fault), .net(N2361), .FEN(FEN[717]), .op(N2361_t2) );
fim FAN_N2361_3 ( .fault(fault), .net(N2361), .FEN(FEN[718]), .op(N2361_t3) );
fim FAN_N2361_4 ( .fault(fault), .net(N2361), .FEN(FEN[719]), .op(N2361_t4) );
fim FAN_N2361_5 ( .fault(fault), .net(N2361), .FEN(FEN[720]), .op(N2361_t5) );
fim FAN_N2361_6 ( .fault(fault), .net(N2361), .FEN(FEN[721]), .op(N2361_t6) );
fim FAN_N2361_7 ( .fault(fault), .net(N2361), .FEN(FEN[722]), .op(N2361_t7) );
fim FAN_N2361_8 ( .fault(fault), .net(N2361), .FEN(FEN[723]), .op(N2361_t8) );
fim FAN_N2361_9 ( .fault(fault), .net(N2361), .FEN(FEN[724]), .op(N2361_t9) );
fim FAN_N2361_10 ( .fault(fault), .net(N2361), .FEN(FEN[725]), .op(N2361_t10) );
fim FAN_N2361_11 ( .fault(fault), .net(N2361), .FEN(FEN[726]), .op(N2361_t11) );
fim FAN_N2361_12 ( .fault(fault), .net(N2361), .FEN(FEN[727]), .op(N2361_t12) );
fim FAN_N2104_0 ( .fault(fault), .net(N2104), .FEN(FEN[728]), .op(N2104_t0) );
fim FAN_N2104_1 ( .fault(fault), .net(N2104), .FEN(FEN[729]), .op(N2104_t1) );
fim FAN_N2104_2 ( .fault(fault), .net(N2104), .FEN(FEN[730]), .op(N2104_t2) );
fim FAN_N2104_3 ( .fault(fault), .net(N2104), .FEN(FEN[731]), .op(N2104_t3) );
fim FAN_N2104_4 ( .fault(fault), .net(N2104), .FEN(FEN[732]), .op(N2104_t4) );
fim FAN_N2104_5 ( .fault(fault), .net(N2104), .FEN(FEN[733]), .op(N2104_t5) );
fim FAN_N2104_6 ( .fault(fault), .net(N2104), .FEN(FEN[734]), .op(N2104_t6) );
fim FAN_N2104_7 ( .fault(fault), .net(N2104), .FEN(FEN[735]), .op(N2104_t7) );
fim FAN_N2104_8 ( .fault(fault), .net(N2104), .FEN(FEN[736]), .op(N2104_t8) );
fim FAN_N2104_9 ( .fault(fault), .net(N2104), .FEN(FEN[737]), .op(N2104_t9) );
fim FAN_N2104_10 ( .fault(fault), .net(N2104), .FEN(FEN[738]), .op(N2104_t10) );
fim FAN_N2104_11 ( .fault(fault), .net(N2104), .FEN(FEN[739]), .op(N2104_t11) );
fim FAN_N2104_12 ( .fault(fault), .net(N2104), .FEN(FEN[740]), .op(N2104_t12) );
fim FAN_N2104_13 ( .fault(fault), .net(N2104), .FEN(FEN[741]), .op(N2104_t13) );
fim FAN_N1171_0 ( .fault(fault), .net(N1171), .FEN(FEN[742]), .op(N1171_t0) );
fim FAN_N1171_1 ( .fault(fault), .net(N1171), .FEN(FEN[743]), .op(N1171_t1) );
fim FAN_N1171_2 ( .fault(fault), .net(N1171), .FEN(FEN[744]), .op(N1171_t2) );
fim FAN_N1171_3 ( .fault(fault), .net(N1171), .FEN(FEN[745]), .op(N1171_t3) );
fim FAN_N1171_4 ( .fault(fault), .net(N1171), .FEN(FEN[746]), .op(N1171_t4) );
fim FAN_N1171_5 ( .fault(fault), .net(N1171), .FEN(FEN[747]), .op(N1171_t5) );
fim FAN_N1171_6 ( .fault(fault), .net(N1171), .FEN(FEN[748]), .op(N1171_t6) );
fim FAN_N1171_7 ( .fault(fault), .net(N1171), .FEN(FEN[749]), .op(N1171_t7) );
fim FAN_N1171_8 ( .fault(fault), .net(N1171), .FEN(FEN[750]), .op(N1171_t8) );
fim FAN_N1171_9 ( .fault(fault), .net(N1171), .FEN(FEN[751]), .op(N1171_t9) );
fim FAN_N1171_10 ( .fault(fault), .net(N1171), .FEN(FEN[752]), .op(N1171_t10) );
fim FAN_N1171_11 ( .fault(fault), .net(N1171), .FEN(FEN[753]), .op(N1171_t11) );
fim FAN_N1171_12 ( .fault(fault), .net(N1171), .FEN(FEN[754]), .op(N1171_t12) );
fim FAN_N1171_13 ( .fault(fault), .net(N1171), .FEN(FEN[755]), .op(N1171_t13) );
fim FAN_N1171_14 ( .fault(fault), .net(N1171), .FEN(FEN[756]), .op(N1171_t14) );
fim FAN_N1171_15 ( .fault(fault), .net(N1171), .FEN(FEN[757]), .op(N1171_t15) );
fim FAN_N2340_0 ( .fault(fault), .net(N2340), .FEN(FEN[758]), .op(N2340_t0) );
fim FAN_N2340_1 ( .fault(fault), .net(N2340), .FEN(FEN[759]), .op(N2340_t1) );
fim FAN_N2340_2 ( .fault(fault), .net(N2340), .FEN(FEN[760]), .op(N2340_t2) );
fim FAN_N2340_3 ( .fault(fault), .net(N2340), .FEN(FEN[761]), .op(N2340_t3) );
fim FAN_N2340_4 ( .fault(fault), .net(N2340), .FEN(FEN[762]), .op(N2340_t4) );
fim FAN_N2340_5 ( .fault(fault), .net(N2340), .FEN(FEN[763]), .op(N2340_t5) );
fim FAN_N2340_6 ( .fault(fault), .net(N2340), .FEN(FEN[764]), .op(N2340_t6) );
fim FAN_N2340_7 ( .fault(fault), .net(N2340), .FEN(FEN[765]), .op(N2340_t7) );
fim FAN_N2340_8 ( .fault(fault), .net(N2340), .FEN(FEN[766]), .op(N2340_t8) );
fim FAN_N2340_9 ( .fault(fault), .net(N2340), .FEN(FEN[767]), .op(N2340_t9) );
fim FAN_N2340_10 ( .fault(fault), .net(N2340), .FEN(FEN[768]), .op(N2340_t10) );
fim FAN_N2340_11 ( .fault(fault), .net(N2340), .FEN(FEN[769]), .op(N2340_t11) );
fim FAN_N2129_0 ( .fault(fault), .net(N2129), .FEN(FEN[770]), .op(N2129_t0) );
fim FAN_N2129_1 ( .fault(fault), .net(N2129), .FEN(FEN[771]), .op(N2129_t1) );
fim FAN_N2129_2 ( .fault(fault), .net(N2129), .FEN(FEN[772]), .op(N2129_t2) );
fim FAN_N2129_3 ( .fault(fault), .net(N2129), .FEN(FEN[773]), .op(N2129_t3) );
fim FAN_N2129_4 ( .fault(fault), .net(N2129), .FEN(FEN[774]), .op(N2129_t4) );
fim FAN_N2129_5 ( .fault(fault), .net(N2129), .FEN(FEN[775]), .op(N2129_t5) );
fim FAN_N2129_6 ( .fault(fault), .net(N2129), .FEN(FEN[776]), .op(N2129_t6) );
fim FAN_N2129_7 ( .fault(fault), .net(N2129), .FEN(FEN[777]), .op(N2129_t7) );
fim FAN_N2129_8 ( .fault(fault), .net(N2129), .FEN(FEN[778]), .op(N2129_t8) );
fim FAN_N2129_9 ( .fault(fault), .net(N2129), .FEN(FEN[779]), .op(N2129_t9) );
fim FAN_N2129_10 ( .fault(fault), .net(N2129), .FEN(FEN[780]), .op(N2129_t10) );
fim FAN_N2129_11 ( .fault(fault), .net(N2129), .FEN(FEN[781]), .op(N2129_t11) );
fim FAN_N2129_12 ( .fault(fault), .net(N2129), .FEN(FEN[782]), .op(N2129_t12) );
fim FAN_N2119_0 ( .fault(fault), .net(N2119), .FEN(FEN[783]), .op(N2119_t0) );
fim FAN_N2119_1 ( .fault(fault), .net(N2119), .FEN(FEN[784]), .op(N2119_t1) );
fim FAN_N2119_2 ( .fault(fault), .net(N2119), .FEN(FEN[785]), .op(N2119_t2) );
fim FAN_N2119_3 ( .fault(fault), .net(N2119), .FEN(FEN[786]), .op(N2119_t3) );
fim FAN_N2119_4 ( .fault(fault), .net(N2119), .FEN(FEN[787]), .op(N2119_t4) );
fim FAN_N2119_5 ( .fault(fault), .net(N2119), .FEN(FEN[788]), .op(N2119_t5) );
fim FAN_N2119_6 ( .fault(fault), .net(N2119), .FEN(FEN[789]), .op(N2119_t6) );
fim FAN_N2119_7 ( .fault(fault), .net(N2119), .FEN(FEN[790]), .op(N2119_t7) );
fim FAN_N2119_8 ( .fault(fault), .net(N2119), .FEN(FEN[791]), .op(N2119_t8) );
fim FAN_N2353_0 ( .fault(fault), .net(N2353), .FEN(FEN[792]), .op(N2353_t0) );
fim FAN_N2353_1 ( .fault(fault), .net(N2353), .FEN(FEN[793]), .op(N2353_t1) );
fim FAN_N2353_2 ( .fault(fault), .net(N2353), .FEN(FEN[794]), .op(N2353_t2) );
fim FAN_N2353_3 ( .fault(fault), .net(N2353), .FEN(FEN[795]), .op(N2353_t3) );
fim FAN_N2353_4 ( .fault(fault), .net(N2353), .FEN(FEN[796]), .op(N2353_t4) );
fim FAN_N2353_5 ( .fault(fault), .net(N2353), .FEN(FEN[797]), .op(N2353_t5) );
fim FAN_N2353_6 ( .fault(fault), .net(N2353), .FEN(FEN[798]), .op(N2353_t6) );
fim FAN_N2297_0 ( .fault(fault), .net(N2297), .FEN(FEN[799]), .op(N2297_t0) );
fim FAN_N2297_1 ( .fault(fault), .net(N2297), .FEN(FEN[800]), .op(N2297_t1) );
fim FAN_N2297_2 ( .fault(fault), .net(N2297), .FEN(FEN[801]), .op(N2297_t2) );
fim FAN_N2297_3 ( .fault(fault), .net(N2297), .FEN(FEN[802]), .op(N2297_t3) );
fim FAN_N2297_4 ( .fault(fault), .net(N2297), .FEN(FEN[803]), .op(N2297_t4) );
fim FAN_N2297_5 ( .fault(fault), .net(N2297), .FEN(FEN[804]), .op(N2297_t5) );
fim FAN_N2297_6 ( .fault(fault), .net(N2297), .FEN(FEN[805]), .op(N2297_t6) );
fim FAN_N2297_7 ( .fault(fault), .net(N2297), .FEN(FEN[806]), .op(N2297_t7) );
fim FAN_N2297_8 ( .fault(fault), .net(N2297), .FEN(FEN[807]), .op(N2297_t8) );
fim FAN_N2297_9 ( .fault(fault), .net(N2297), .FEN(FEN[808]), .op(N2297_t9) );
fim FAN_N2297_10 ( .fault(fault), .net(N2297), .FEN(FEN[809]), .op(N2297_t10) );
fim FAN_N2297_11 ( .fault(fault), .net(N2297), .FEN(FEN[810]), .op(N2297_t11) );
fim FAN_N2297_12 ( .fault(fault), .net(N2297), .FEN(FEN[811]), .op(N2297_t12) );
fim FAN_N2297_13 ( .fault(fault), .net(N2297), .FEN(FEN[812]), .op(N2297_t13) );
fim FAN_N2297_14 ( .fault(fault), .net(N2297), .FEN(FEN[813]), .op(N2297_t14) );
fim FAN_N2375_0 ( .fault(fault), .net(N2375), .FEN(FEN[814]), .op(N2375_t0) );
fim FAN_N2375_1 ( .fault(fault), .net(N2375), .FEN(FEN[815]), .op(N2375_t1) );
fim FAN_N2375_2 ( .fault(fault), .net(N2375), .FEN(FEN[816]), .op(N2375_t2) );
fim FAN_N2375_3 ( .fault(fault), .net(N2375), .FEN(FEN[817]), .op(N2375_t3) );
fim FAN_N2375_4 ( .fault(fault), .net(N2375), .FEN(FEN[818]), .op(N2375_t4) );
fim FAN_N2375_5 ( .fault(fault), .net(N2375), .FEN(FEN[819]), .op(N2375_t5) );
fim FAN_N2375_6 ( .fault(fault), .net(N2375), .FEN(FEN[820]), .op(N2375_t6) );
fim FAN_N2375_7 ( .fault(fault), .net(N2375), .FEN(FEN[821]), .op(N2375_t7) );
fim FAN_N1188_0 ( .fault(fault), .net(N1188), .FEN(FEN[822]), .op(N1188_t0) );
fim FAN_N1188_1 ( .fault(fault), .net(N1188), .FEN(FEN[823]), .op(N1188_t1) );
fim FAN_N1188_2 ( .fault(fault), .net(N1188), .FEN(FEN[824]), .op(N1188_t2) );
fim FAN_N1188_3 ( .fault(fault), .net(N1188), .FEN(FEN[825]), .op(N1188_t3) );
fim FAN_N1188_4 ( .fault(fault), .net(N1188), .FEN(FEN[826]), .op(N1188_t4) );
fim FAN_N1188_5 ( .fault(fault), .net(N1188), .FEN(FEN[827]), .op(N1188_t5) );
fim FAN_N1188_6 ( .fault(fault), .net(N1188), .FEN(FEN[828]), .op(N1188_t6) );
fim FAN_N1188_7 ( .fault(fault), .net(N1188), .FEN(FEN[829]), .op(N1188_t7) );
fim FAN_N1188_8 ( .fault(fault), .net(N1188), .FEN(FEN[830]), .op(N1188_t8) );
fim FAN_N1188_9 ( .fault(fault), .net(N1188), .FEN(FEN[831]), .op(N1188_t9) );
fim FAN_N1188_10 ( .fault(fault), .net(N1188), .FEN(FEN[832]), .op(N1188_t10) );
fim FAN_N1188_11 ( .fault(fault), .net(N1188), .FEN(FEN[833]), .op(N1188_t11) );
fim FAN_N1188_12 ( .fault(fault), .net(N1188), .FEN(FEN[834]), .op(N1188_t12) );
fim FAN_N1188_13 ( .fault(fault), .net(N1188), .FEN(FEN[835]), .op(N1188_t13) );
fim FAN_N1188_14 ( .fault(fault), .net(N1188), .FEN(FEN[836]), .op(N1188_t14) );
fim FAN_N1188_15 ( .fault(fault), .net(N1188), .FEN(FEN[837]), .op(N1188_t15) );
fim FAN_N2326_0 ( .fault(fault), .net(N2326), .FEN(FEN[838]), .op(N2326_t0) );
fim FAN_N2326_1 ( .fault(fault), .net(N2326), .FEN(FEN[839]), .op(N2326_t1) );
fim FAN_N2326_2 ( .fault(fault), .net(N2326), .FEN(FEN[840]), .op(N2326_t2) );
fim FAN_N2326_3 ( .fault(fault), .net(N2326), .FEN(FEN[841]), .op(N2326_t3) );
fim FAN_N2326_4 ( .fault(fault), .net(N2326), .FEN(FEN[842]), .op(N2326_t4) );
fim FAN_N2326_5 ( .fault(fault), .net(N2326), .FEN(FEN[843]), .op(N2326_t5) );
fim FAN_N2326_6 ( .fault(fault), .net(N2326), .FEN(FEN[844]), .op(N2326_t6) );
fim FAN_N2326_7 ( .fault(fault), .net(N2326), .FEN(FEN[845]), .op(N2326_t7) );
fim FAN_N2326_8 ( .fault(fault), .net(N2326), .FEN(FEN[846]), .op(N2326_t8) );
fim FAN_N2326_9 ( .fault(fault), .net(N2326), .FEN(FEN[847]), .op(N2326_t9) );
fim FAN_N2326_10 ( .fault(fault), .net(N2326), .FEN(FEN[848]), .op(N2326_t10) );
fim FAN_N2326_11 ( .fault(fault), .net(N2326), .FEN(FEN[849]), .op(N2326_t11) );
fim FAN_N2326_12 ( .fault(fault), .net(N2326), .FEN(FEN[850]), .op(N2326_t12) );
fim FAN_N2143_0 ( .fault(fault), .net(N2143), .FEN(FEN[851]), .op(N2143_t0) );
fim FAN_N2143_1 ( .fault(fault), .net(N2143), .FEN(FEN[852]), .op(N2143_t1) );
fim FAN_N2143_2 ( .fault(fault), .net(N2143), .FEN(FEN[853]), .op(N2143_t2) );
fim FAN_N2143_3 ( .fault(fault), .net(N2143), .FEN(FEN[854]), .op(N2143_t3) );
fim FAN_N2427_0 ( .fault(fault), .net(N2427), .FEN(FEN[855]), .op(N2427_t0) );
fim FAN_N2427_1 ( .fault(fault), .net(N2427), .FEN(FEN[856]), .op(N2427_t1) );
fim FAN_N2427_2 ( .fault(fault), .net(N2427), .FEN(FEN[857]), .op(N2427_t2) );
fim FAN_N2427_3 ( .fault(fault), .net(N2427), .FEN(FEN[858]), .op(N2427_t3) );
fim FAN_N2427_4 ( .fault(fault), .net(N2427), .FEN(FEN[859]), .op(N2427_t4) );
fim FAN_N2427_5 ( .fault(fault), .net(N2427), .FEN(FEN[860]), .op(N2427_t5) );
fim FAN_N2427_6 ( .fault(fault), .net(N2427), .FEN(FEN[861]), .op(N2427_t6) );
fim FAN_N2427_7 ( .fault(fault), .net(N2427), .FEN(FEN[862]), .op(N2427_t7) );
fim FAN_N2427_8 ( .fault(fault), .net(N2427), .FEN(FEN[863]), .op(N2427_t8) );
fim FAN_N2427_9 ( .fault(fault), .net(N2427), .FEN(FEN[864]), .op(N2427_t9) );
fim FAN_N2427_10 ( .fault(fault), .net(N2427), .FEN(FEN[865]), .op(N2427_t10) );
fim FAN_N2427_11 ( .fault(fault), .net(N2427), .FEN(FEN[866]), .op(N2427_t11) );
fim FAN_N2427_12 ( .fault(fault), .net(N2427), .FEN(FEN[867]), .op(N2427_t12) );
fim FAN_N2427_13 ( .fault(fault), .net(N2427), .FEN(FEN[868]), .op(N2427_t13) );
fim FAN_N2427_14 ( .fault(fault), .net(N2427), .FEN(FEN[869]), .op(N2427_t14) );
fim FAN_N2427_15 ( .fault(fault), .net(N2427), .FEN(FEN[870]), .op(N2427_t15) );
fim FAN_N2386_0 ( .fault(fault), .net(N2386), .FEN(FEN[871]), .op(N2386_t0) );
fim FAN_N2386_1 ( .fault(fault), .net(N2386), .FEN(FEN[872]), .op(N2386_t1) );
fim FAN_N2386_2 ( .fault(fault), .net(N2386), .FEN(FEN[873]), .op(N2386_t2) );
fim FAN_N2386_3 ( .fault(fault), .net(N2386), .FEN(FEN[874]), .op(N2386_t3) );
fim FAN_N2386_4 ( .fault(fault), .net(N2386), .FEN(FEN[875]), .op(N2386_t4) );
fim FAN_N2386_5 ( .fault(fault), .net(N2386), .FEN(FEN[876]), .op(N2386_t5) );
fim FAN_N2386_6 ( .fault(fault), .net(N2386), .FEN(FEN[877]), .op(N2386_t6) );
fim FAN_N2386_7 ( .fault(fault), .net(N2386), .FEN(FEN[878]), .op(N2386_t7) );
fim FAN_N2386_8 ( .fault(fault), .net(N2386), .FEN(FEN[879]), .op(N2386_t8) );
fim FAN_N2386_9 ( .fault(fault), .net(N2386), .FEN(FEN[880]), .op(N2386_t9) );
fim FAN_N2386_10 ( .fault(fault), .net(N2386), .FEN(FEN[881]), .op(N2386_t10) );
fim FAN_N2386_11 ( .fault(fault), .net(N2386), .FEN(FEN[882]), .op(N2386_t11) );
fim FAN_N2386_12 ( .fault(fault), .net(N2386), .FEN(FEN[883]), .op(N2386_t12) );
fim FAN_N2386_13 ( .fault(fault), .net(N2386), .FEN(FEN[884]), .op(N2386_t13) );
fim FAN_N926_0 ( .fault(fault), .net(N926), .FEN(FEN[885]), .op(N926_t0) );
fim FAN_N926_1 ( .fault(fault), .net(N926), .FEN(FEN[886]), .op(N926_t1) );
fim FAN_N926_2 ( .fault(fault), .net(N926), .FEN(FEN[887]), .op(N926_t2) );
fim FAN_N926_3 ( .fault(fault), .net(N926), .FEN(FEN[888]), .op(N926_t3) );
fim FAN_N926_4 ( .fault(fault), .net(N926), .FEN(FEN[889]), .op(N926_t4) );
fim FAN_N926_5 ( .fault(fault), .net(N926), .FEN(FEN[890]), .op(N926_t5) );
fim FAN_N926_6 ( .fault(fault), .net(N926), .FEN(FEN[891]), .op(N926_t6) );
fim FAN_N926_7 ( .fault(fault), .net(N926), .FEN(FEN[892]), .op(N926_t7) );
fim FAN_N2558_0 ( .fault(fault), .net(N2558), .FEN(FEN[893]), .op(N2558_t0) );
fim FAN_N2558_1 ( .fault(fault), .net(N2558), .FEN(FEN[894]), .op(N2558_t1) );
fim FAN_N2561_0 ( .fault(fault), .net(N2561), .FEN(FEN[895]), .op(N2561_t0) );
fim FAN_N2561_1 ( .fault(fault), .net(N2561), .FEN(FEN[896]), .op(N2561_t1) );
fim FAN_N2564_0 ( .fault(fault), .net(N2564), .FEN(FEN[897]), .op(N2564_t0) );
fim FAN_N2564_1 ( .fault(fault), .net(N2564), .FEN(FEN[898]), .op(N2564_t1) );
fim FAN_N2567_0 ( .fault(fault), .net(N2567), .FEN(FEN[899]), .op(N2567_t0) );
fim FAN_N2567_1 ( .fault(fault), .net(N2567), .FEN(FEN[900]), .op(N2567_t1) );
fim FAN_N2570_0 ( .fault(fault), .net(N2570), .FEN(FEN[901]), .op(N2570_t0) );
fim FAN_N2570_1 ( .fault(fault), .net(N2570), .FEN(FEN[902]), .op(N2570_t1) );
fim FAN_N2573_0 ( .fault(fault), .net(N2573), .FEN(FEN[903]), .op(N2573_t0) );
fim FAN_N2573_1 ( .fault(fault), .net(N2573), .FEN(FEN[904]), .op(N2573_t1) );
fim FAN_N2576_0 ( .fault(fault), .net(N2576), .FEN(FEN[905]), .op(N2576_t0) );
fim FAN_N2576_1 ( .fault(fault), .net(N2576), .FEN(FEN[906]), .op(N2576_t1) );
fim FAN_N2639_0 ( .fault(fault), .net(N2639), .FEN(FEN[907]), .op(N2639_t0) );
fim FAN_N2639_1 ( .fault(fault), .net(N2639), .FEN(FEN[908]), .op(N2639_t1) );
fim FAN_N2642_0 ( .fault(fault), .net(N2642), .FEN(FEN[909]), .op(N2642_t0) );
fim FAN_N2642_1 ( .fault(fault), .net(N2642), .FEN(FEN[910]), .op(N2642_t1) );
fim FAN_N2645_0 ( .fault(fault), .net(N2645), .FEN(FEN[911]), .op(N2645_t0) );
fim FAN_N2645_1 ( .fault(fault), .net(N2645), .FEN(FEN[912]), .op(N2645_t1) );
fim FAN_N2648_0 ( .fault(fault), .net(N2648), .FEN(FEN[913]), .op(N2648_t0) );
fim FAN_N2648_1 ( .fault(fault), .net(N2648), .FEN(FEN[914]), .op(N2648_t1) );
fim FAN_N2651_0 ( .fault(fault), .net(N2651), .FEN(FEN[915]), .op(N2651_t0) );
fim FAN_N2651_1 ( .fault(fault), .net(N2651), .FEN(FEN[916]), .op(N2651_t1) );
fim FAN_N2655_0 ( .fault(fault), .net(N2655), .FEN(FEN[917]), .op(N2655_t0) );
fim FAN_N2655_1 ( .fault(fault), .net(N2655), .FEN(FEN[918]), .op(N2655_t1) );
fim FAN_N2658_0 ( .fault(fault), .net(N2658), .FEN(FEN[919]), .op(N2658_t0) );
fim FAN_N2658_1 ( .fault(fault), .net(N2658), .FEN(FEN[920]), .op(N2658_t1) );
fim FAN_N2661_0 ( .fault(fault), .net(N2661), .FEN(FEN[921]), .op(N2661_t0) );
fim FAN_N2661_1 ( .fault(fault), .net(N2661), .FEN(FEN[922]), .op(N2661_t1) );
fim FAN_N2664_0 ( .fault(fault), .net(N2664), .FEN(FEN[923]), .op(N2664_t0) );
fim FAN_N2664_1 ( .fault(fault), .net(N2664), .FEN(FEN[924]), .op(N2664_t1) );
fim FAN_N2537_0 ( .fault(fault), .net(N2537), .FEN(FEN[925]), .op(N2537_t0) );
fim FAN_N2537_1 ( .fault(fault), .net(N2537), .FEN(FEN[926]), .op(N2537_t1) );
fim FAN_N2540_0 ( .fault(fault), .net(N2540), .FEN(FEN[927]), .op(N2540_t0) );
fim FAN_N2540_1 ( .fault(fault), .net(N2540), .FEN(FEN[928]), .op(N2540_t1) );
fim FAN_N2543_0 ( .fault(fault), .net(N2543), .FEN(FEN[929]), .op(N2543_t0) );
fim FAN_N2543_1 ( .fault(fault), .net(N2543), .FEN(FEN[930]), .op(N2543_t1) );
fim FAN_N2546_0 ( .fault(fault), .net(N2546), .FEN(FEN[931]), .op(N2546_t0) );
fim FAN_N2546_1 ( .fault(fault), .net(N2546), .FEN(FEN[932]), .op(N2546_t1) );
fim FAN_N2594_0 ( .fault(fault), .net(N2594), .FEN(FEN[933]), .op(N2594_t0) );
fim FAN_N2594_1 ( .fault(fault), .net(N2594), .FEN(FEN[934]), .op(N2594_t1) );
fim FAN_N2597_0 ( .fault(fault), .net(N2597), .FEN(FEN[935]), .op(N2597_t0) );
fim FAN_N2597_1 ( .fault(fault), .net(N2597), .FEN(FEN[936]), .op(N2597_t1) );
fim FAN_N2600_0 ( .fault(fault), .net(N2600), .FEN(FEN[937]), .op(N2600_t0) );
fim FAN_N2600_1 ( .fault(fault), .net(N2600), .FEN(FEN[938]), .op(N2600_t1) );
fim FAN_N2603_0 ( .fault(fault), .net(N2603), .FEN(FEN[939]), .op(N2603_t0) );
fim FAN_N2603_1 ( .fault(fault), .net(N2603), .FEN(FEN[940]), .op(N2603_t1) );
fim FAN_N2606_0 ( .fault(fault), .net(N2606), .FEN(FEN[941]), .op(N2606_t0) );
fim FAN_N2606_1 ( .fault(fault), .net(N2606), .FEN(FEN[942]), .op(N2606_t1) );
fim FAN_N2549_0 ( .fault(fault), .net(N2549), .FEN(FEN[943]), .op(N2549_t0) );
fim FAN_N2549_1 ( .fault(fault), .net(N2549), .FEN(FEN[944]), .op(N2549_t1) );
fim FAN_N2611_0 ( .fault(fault), .net(N2611), .FEN(FEN[945]), .op(N2611_t0) );
fim FAN_N2611_1 ( .fault(fault), .net(N2611), .FEN(FEN[946]), .op(N2611_t1) );
fim FAN_N2614_0 ( .fault(fault), .net(N2614), .FEN(FEN[947]), .op(N2614_t0) );
fim FAN_N2614_1 ( .fault(fault), .net(N2614), .FEN(FEN[948]), .op(N2614_t1) );
fim FAN_N2617_0 ( .fault(fault), .net(N2617), .FEN(FEN[949]), .op(N2617_t0) );
fim FAN_N2617_1 ( .fault(fault), .net(N2617), .FEN(FEN[950]), .op(N2617_t1) );
fim FAN_N2620_0 ( .fault(fault), .net(N2620), .FEN(FEN[951]), .op(N2620_t0) );
fim FAN_N2620_1 ( .fault(fault), .net(N2620), .FEN(FEN[952]), .op(N2620_t1) );
fim FAN_N2552_0 ( .fault(fault), .net(N2552), .FEN(FEN[953]), .op(N2552_t0) );
fim FAN_N2552_1 ( .fault(fault), .net(N2552), .FEN(FEN[954]), .op(N2552_t1) );
fim FAN_N2555_0 ( .fault(fault), .net(N2555), .FEN(FEN[955]), .op(N2555_t0) );
fim FAN_N2555_1 ( .fault(fault), .net(N2555), .FEN(FEN[956]), .op(N2555_t1) );
fim FAN_N2747_0 ( .fault(fault), .net(N2747), .FEN(FEN[957]), .op(N2747_t0) );
fim FAN_N2747_1 ( .fault(fault), .net(N2747), .FEN(FEN[958]), .op(N2747_t1) );
fim FAN_N2750_0 ( .fault(fault), .net(N2750), .FEN(FEN[959]), .op(N2750_t0) );
fim FAN_N2750_1 ( .fault(fault), .net(N2750), .FEN(FEN[960]), .op(N2750_t1) );
fim FAN_N2773_0 ( .fault(fault), .net(N2773), .FEN(FEN[961]), .op(N2773_t0) );
fim FAN_N2773_1 ( .fault(fault), .net(N2773), .FEN(FEN[962]), .op(N2773_t1) );
fim FAN_N2776_0 ( .fault(fault), .net(N2776), .FEN(FEN[963]), .op(N2776_t0) );
fim FAN_N2776_1 ( .fault(fault), .net(N2776), .FEN(FEN[964]), .op(N2776_t1) );
fim FAN_N283_0 ( .fault(fault), .net(N283), .FEN(FEN[965]), .op(N283_t0) );
fim FAN_N283_1 ( .fault(fault), .net(N283), .FEN(FEN[966]), .op(N283_t1) );
fim FAN_N283_2 ( .fault(fault), .net(N283), .FEN(FEN[967]), .op(N283_t2) );
fim FAN_N283_3 ( .fault(fault), .net(N283), .FEN(FEN[968]), .op(N283_t3) );
fim FAN_N283_4 ( .fault(fault), .net(N283), .FEN(FEN[969]), .op(N283_t4) );
fim FAN_N283_5 ( .fault(fault), .net(N283), .FEN(FEN[970]), .op(N283_t5) );
fim FAN_N2789_0 ( .fault(fault), .net(N2789), .FEN(FEN[971]), .op(N2789_t0) );
fim FAN_N2789_1 ( .fault(fault), .net(N2789), .FEN(FEN[972]), .op(N2789_t1) );
fim FAN_N2789_2 ( .fault(fault), .net(N2789), .FEN(FEN[973]), .op(N2789_t2) );
fim FAN_N2789_3 ( .fault(fault), .net(N2789), .FEN(FEN[974]), .op(N2789_t3) );
fim FAN_N2789_4 ( .fault(fault), .net(N2789), .FEN(FEN[975]), .op(N2789_t4) );
fim FAN_N2789_5 ( .fault(fault), .net(N2789), .FEN(FEN[976]), .op(N2789_t5) );
fim FAN_N2812_0 ( .fault(fault), .net(N2812), .FEN(FEN[977]), .op(N2812_t0) );
fim FAN_N2812_1 ( .fault(fault), .net(N2812), .FEN(FEN[978]), .op(N2812_t1) );
fim FAN_N2815_0 ( .fault(fault), .net(N2815), .FEN(FEN[979]), .op(N2815_t0) );
fim FAN_N2815_1 ( .fault(fault), .net(N2815), .FEN(FEN[980]), .op(N2815_t1) );
fim FAN_N2818_0 ( .fault(fault), .net(N2818), .FEN(FEN[981]), .op(N2818_t0) );
fim FAN_N2818_1 ( .fault(fault), .net(N2818), .FEN(FEN[982]), .op(N2818_t1) );
fim FAN_N2821_0 ( .fault(fault), .net(N2821), .FEN(FEN[983]), .op(N2821_t0) );
fim FAN_N2821_1 ( .fault(fault), .net(N2821), .FEN(FEN[984]), .op(N2821_t1) );
fim FAN_N2824_0 ( .fault(fault), .net(N2824), .FEN(FEN[985]), .op(N2824_t0) );
fim FAN_N2824_1 ( .fault(fault), .net(N2824), .FEN(FEN[986]), .op(N2824_t1) );
fim FAN_N2829_0 ( .fault(fault), .net(N2829), .FEN(FEN[987]), .op(N2829_t0) );
fim FAN_N2829_1 ( .fault(fault), .net(N2829), .FEN(FEN[988]), .op(N2829_t1) );
fim FAN_N2843_0 ( .fault(fault), .net(N2843), .FEN(FEN[989]), .op(N2843_t0) );
fim FAN_N2843_1 ( .fault(fault), .net(N2843), .FEN(FEN[990]), .op(N2843_t1) );
fim FAN_N2846_0 ( .fault(fault), .net(N2846), .FEN(FEN[991]), .op(N2846_t0) );
fim FAN_N2846_1 ( .fault(fault), .net(N2846), .FEN(FEN[992]), .op(N2846_t1) );
fim FAN_N2883_0 ( .fault(fault), .net(N2883), .FEN(FEN[993]), .op(N2883_t0) );
fim FAN_N2883_1 ( .fault(fault), .net(N2883), .FEN(FEN[994]), .op(N2883_t1) );
initial begin
    FEN <= {994'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {994'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,994'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,994'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN = {FEN[993:0], FEN[994]};
        if( ((FEN[361] || FEN[364]) && fault == 0) || ((FEN[221] || FEN[224] || FEN[250] || FEN[252] || FEN[689]) && fault)) FEN = {FEN[993:0], FEN[994]};
        if (FEN[690] && fault) FEN = {FEN[993:0], FEN[994]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
    // EndFaultModel

//Anchor
not NOT1_1 (N190, N1_t0);
not NOT1_2 (N194, N4_t0);
not NOT1_3 (N197, N7_t0);
not NOT1_4 (N201, N10_t0);
not NOT1_5 (N206, N13_t0);
not NOT1_6 (N209, N16_t0);
not NOT1_7 (N212, N19_t0);
not NOT1_8 (N216, N22_t0);
not NOT1_9 (N220, N25_t0);
not NOT1_10 (N225, N28_t0);
not NOT1_11 (N229, N31_t0);
not NOT1_12 (N232, N34_t0);
not NOT1_13 (N235, N37_t0);
not NOT1_14 (N239, N40_t0);
not NOT1_15 (N243, N43_t0);
not NOT1_16 (N247, N46_t0);
nand NAND2_17 (N251, N63_t0, N88_t0);
nand NAND2_18 (N252, N66_t0, N91_t0);
not NOT1_19 (N253, N72_t0);
not NOT1_20 (N256, N72_t1);
buf BUFF1_21 (N257, N69_t0);
buf BUFF1_22 (N260, N69_t1);
not NOT1_23 (N263, N76_t0);
not NOT1_24 (N266, N79_t0);
not NOT1_25 (N269, N82_t0);
not NOT1_26 (N272, N85_t0);
not NOT1_27 (N275, N104_t0);
not NOT1_28 (N276, N104_t1);
not NOT1_29 (N277, N88_t1);
not NOT1_30 (N280, N91_t1);
buf BUFF1_31 (N283, N94_t0);
not NOT1_32 (N290, N94_t1);
buf BUFF1_33 (N297, N94_t2);
not NOT1_34 (N300, N94_t3);
buf BUFF1_35 (N303, N99_t0);
not NOT1_36 (N306, N99_t1);
not NOT1_37 (N313, N99_t2);
buf BUFF1_38 (N316, N104_t2);
not NOT1_39 (N319, N104_t3);
buf BUFF1_40 (N326, N104_t4);
buf BUFF1_41 (N331, N104_t5);
not NOT1_42 (N338, N104_t6);
buf BUFF1_43 (N343, N1_t1);
buf BUFF1_44 (N346, N4_t1);
buf BUFF1_45 (N349, N7_t1);
buf BUFF1_46 (N352, N10_t1);
buf BUFF1_47 (N355, N13_t1);
buf BUFF1_48 (N358, N16_t1);
buf BUFF1_49 (N361, N19_t1);
buf BUFF1_50 (N364, N22_t1);
buf BUFF1_51 (N367, N25_t1);
buf BUFF1_52 (N370, N28_t1);
buf BUFF1_53 (N373, N31_t1);
buf BUFF1_54 (N376, N34_t1);
buf BUFF1_55 (N379, N37_t1);
buf BUFF1_56 (N382, N40_t1);
buf BUFF1_57 (N385, N43_t1);
buf BUFF1_58 (N388, N46_t1);
not NOT1_59 (N534, N343_t0);
not NOT1_60 (N535, N346_t0);
not NOT1_61 (N536, N349_t0);
not NOT1_62 (N537, N352_t0);
not NOT1_63 (N538, N355_t0);
not NOT1_64 (N539, N358_t0);
not NOT1_65 (N540, N361_t0);
not NOT1_66 (N541, N364_t0);
not NOT1_67 (N542, N367_t0);
not NOT1_68 (N543, N370_t0);
not NOT1_69 (N544, N373_t0);
not NOT1_70 (N545, N376_t0);
not NOT1_71 (N546, N379_t0);
not NOT1_72 (N547, N382_t0);
not NOT1_73 (N548, N385_t0);
not NOT1_74 (N549, N388_t0);
nand NAND2_75 (N550, N306_t0, N331_t0);
nand NAND2_76 (N551, N306_t1, N331_t1);
nand NAND2_77 (N552, N306_t2, N331_t2);
nand NAND2_78 (N553, N306_t3, N331_t3);
nand NAND2_79 (N554, N306_t4, N331_t4);
nand NAND2_80 (N555, N306_t5, N331_t5);
buf BUFF1_81 (N556, N190_t0);
buf BUFF1_82 (N559, N194_t0);
buf BUFF1_83 (N562, N206_t0);
buf BUFF1_84 (N565, N209_t0);
buf BUFF1_85 (N568, N225_t0);
buf BUFF1_86 (N571, N243_t0);
and AND2_87 (N574, N63_t1, N319_t0);
buf BUFF1_88 (N577, N220_t0);
buf BUFF1_89 (N580, N229_t0);
buf BUFF1_90 (N583, N232_t0);
and AND2_91 (N586, N66_t1, N319_t1);
buf BUFF1_92 (N589, N239_t0);
and AND3_93 (N592, N49_t0, N253_t0, N319_t2);
buf BUFF1_94 (N595, N247_t0);
buf BUFF1_95 (N598, N239_t1);
nand NAND2_96 (N601, N326_t0, N277_t0);
nand NAND2_97 (N602, N326_t1, N280_t0);
nand NAND2_98 (N603, N260_t0, N72_t2);
nand NAND2_99 (N608, N260_t1, N300_t0);
nand NAND2_100 (N612, N256, N300_t1);
buf BUFF1_101 (N616, N201_t0);
buf BUFF1_102 (N619, N216_t0);
buf BUFF1_103 (N622, N220_t1);
buf BUFF1_104 (N625, N239_t2);
buf BUFF1_105 (N628, N190_t1);
buf BUFF1_106 (N631, N190_t2);
buf BUFF1_107 (N634, N194_t1);
buf BUFF1_108 (N637, N229_t1);
buf BUFF1_109 (N640, N197_t0);
and AND3_110 (N643, N56_t0, N257_t0, N319_t3);
buf BUFF1_111 (N646, N232_t1);
buf BUFF1_112 (N649, N201_t1);
buf BUFF1_113 (N652, N235_t0);
and AND3_114 (N655, N60_t0, N257_t1, N319_t4);
buf BUFF1_115 (N658, N263_t0);
buf BUFF1_116 (N661, N263_t1);
buf BUFF1_117 (N664, N266_t0);
buf BUFF1_118 (N667, N266_t1);
buf BUFF1_119 (N670, N269_t0);
buf BUFF1_120 (N673, N269_t1);
buf BUFF1_121 (N676, N272_t0);
buf BUFF1_122 (N679, N272_t1);
and AND2_123 (N682, N251, N316_t0);
and AND2_124 (N685, N252, N316_t1);
buf BUFF1_125 (N688, N197_t1);
buf BUFF1_126 (N691, N197_t2);
buf BUFF1_127 (N694, N212_t0);
buf BUFF1_128 (N697, N212_t1);
buf BUFF1_129 (N700, N247_t1);
buf BUFF1_130 (N703, N247_t2);
buf BUFF1_131 (N706, N235_t1);
buf BUFF1_132 (N709, N235_t2);
buf BUFF1_133 (N712, N201_t2);
buf BUFF1_134 (N715, N201_t3);
buf BUFF1_135 (N718, N206_t1);
buf BUFF1_136 (N721, N216_t1);
and AND3_137 (N724, N53_t0, N253_t1, N319_t5);
buf BUFF1_138 (N727, N243_t1);
buf BUFF1_139 (N730, N220_t2);
buf BUFF1_140 (N733, N220_t3);
buf BUFF1_141 (N736, N209_t1);
buf BUFF1_142 (N739, N216_t2);
buf BUFF1_143 (N742, N225_t1);
buf BUFF1_144 (N745, N243_t2);
buf BUFF1_145 (N748, N212_t2);
buf BUFF1_146 (N751, N225_t2);
not NOT1_147 (N886, N682_t0);
not NOT1_148 (N887, N685_t0);
not NOT1_149 (N888, N616_t0);
not NOT1_150 (N889, N619_t0);
not NOT1_151 (N890, N622_t0);
not NOT1_152 (N891, N625_t0);
not NOT1_153 (N892, N631_t0);
not NOT1_154 (N893, N643_t0);
not NOT1_155 (N894, N649_t0);
not NOT1_156 (N895, N652_t0);
not NOT1_157 (N896, N655_t0);
and AND2_158 (N897, N49_t1, N612_t0);
and AND2_159 (N898, N56_t1, N608_t0);
nand NAND2_160 (N899, N53_t1, N612_t1);
nand NAND2_161 (N903, N60_t1, N608_t1);
nand NAND2_162 (N907, N49_t2, N612_t2);
nand NAND2_163 (N910, N56_t2, N608_t2);
not NOT1_164 (N913, N661_t0);
not NOT1_165 (N914, N658_t0);
not NOT1_166 (N915, N667_t0);
not NOT1_167 (N916, N664_t0);
not NOT1_168 (N917, N673_t0);
not NOT1_169 (N918, N670_t0);
not NOT1_170 (N919, N679_t0);
not NOT1_171 (N920, N676_t0);
nand NAND4_172 (N921, N277_t1, N297_t0, N326_t2, N603_t0);
nand NAND4_173 (N922, N280_t1, N297_t1, N326_t3, N603_t1);
nand NAND3_174 (N923, N303_t0, N338_t0, N603_t2);
and AND3_175 (N926, N303_t1, N338_t1, N603_t3);
buf BUFF1_176 (N935, N556_t0);
not NOT1_177 (N938, N688_t0);
buf BUFF1_178 (N939, N556_t1);
not NOT1_179 (N942, N691_t0);
buf BUFF1_180 (N943, N562_t0);
not NOT1_181 (N946, N694_t0);
buf BUFF1_182 (N947, N562_t1);
not NOT1_183 (N950, N697_t0);
buf BUFF1_184 (N951, N568_t0);
not NOT1_185 (N954, N700_t0);
buf BUFF1_186 (N955, N568_t1);
not NOT1_187 (N958, N703_t0);
buf BUFF1_188 (N959, N574_t0);
buf BUFF1_189 (N962, N574_t1);
buf BUFF1_190 (N965, N580_t0);
not NOT1_191 (N968, N706_t0);
buf BUFF1_192 (N969, N580_t1);
not NOT1_193 (N972, N709_t0);
buf BUFF1_194 (N973, N586_t0);
not NOT1_195 (N976, N712_t0);
buf BUFF1_196 (N977, N586_t1);
not NOT1_197 (N980, N715_t0);
buf BUFF1_198 (N981, N592_t0);
not NOT1_199 (N984, N628_t0);
buf BUFF1_200 (N985, N592_t1);
not NOT1_201 (N988, N718_t0);
not NOT1_202 (N989, N721_t0);
not NOT1_203 (N990, N634_t0);
not NOT1_204 (N991, N724_t0);
not NOT1_205 (N992, N727_t0);
not NOT1_206 (N993, N637_t0);
buf BUFF1_207 (N994, N595_t0);
not NOT1_208 (N997, N730_t0);
buf BUFF1_209 (N998, N595_t1);
not NOT1_210 (N1001, N733_t0);
not NOT1_211 (N1002, N736_t0);
not NOT1_212 (N1003, N739_t0);
not NOT1_213 (N1004, N640_t0);
not NOT1_214 (N1005, N742_t0);
not NOT1_215 (N1006, N745_t0);
not NOT1_216 (N1007, N646_t0);
not NOT1_217 (N1008, N748_t0);
not NOT1_218 (N1009, N751_t0);
buf BUFF1_219 (N1010, N559_t0);
buf BUFF1_220 (N1013, N559_t1);
buf BUFF1_221 (N1016, N565_t0);
buf BUFF1_222 (N1019, N565_t1);
buf BUFF1_223 (N1022, N571_t0);
buf BUFF1_224 (N1025, N571_t1);
buf BUFF1_225 (N1028, N577_t0);
buf BUFF1_226 (N1031, N577_t1);
buf BUFF1_227 (N1034, N583_t0);
buf BUFF1_228 (N1037, N583_t1);
buf BUFF1_229 (N1040, N589_t0);
buf BUFF1_230 (N1043, N589_t1);
buf BUFF1_231 (N1046, N598_t0);
buf BUFF1_232 (N1049, N598_t1);
nand NAND2_233 (N1054, N619_t1, N888);
nand NAND2_234 (N1055, N616_t1, N889);
nand NAND2_235 (N1063, N625_t1, N890);
nand NAND2_236 (N1064, N622_t1, N891);
nand NAND2_237 (N1067, N655_t1, N895);
nand NAND2_238 (N1068, N652_t1, N896);
nand NAND2_239 (N1119, N721_t1, N988);
nand NAND2_240 (N1120, N718_t1, N989);
nand NAND2_241 (N1121, N727_t1, N991);
nand NAND2_242 (N1122, N724_t1, N992);
nand NAND2_243 (N1128, N739_t1, N1002);
nand NAND2_244 (N1129, N736_t1, N1003);
nand NAND2_245 (N1130, N745_t1, N1005);
nand NAND2_246 (N1131, N742_t1, N1006);
nand NAND2_247 (N1132, N751_t1, N1008);
nand NAND2_248 (N1133, N748_t1, N1009);
not NOT1_249 (N1148, N939_t0);
not NOT1_250 (N1149, N935_t0);
nand NAND2_251 (N1150, N1054, N1055);
not NOT1_252 (N1151, N943_t0);
not NOT1_253 (N1152, N947_t0);
not NOT1_254 (N1153, N955_t0);
not NOT1_255 (N1154, N951_t0);
not NOT1_256 (N1155, N962_t0);
not NOT1_257 (N1156, N969_t0);
not NOT1_258 (N1157, N977_t0);
nand NAND2_259 (N1158, N1063, N1064);
not NOT1_260 (N1159, N985_t0);
nand NAND2_261 (N1160, N985_t1, N892);
not NOT1_262 (N1161, N998_t0);
nand NAND2_263 (N1162, N1067, N1068);
not NOT1_264 (N1163, N899_t0);
buf BUFF1_265 (N1164, N899_t1);
not NOT1_266 (N1167, N903_t0);
buf BUFF1_267 (N1168, N903_t1);
nand NAND2_268 (N1171, N921, N923_t0);
nand NAND2_269 (N1188, N922, N923_t1);
not NOT1_270 (N1205, N1010_t0);
nand NAND2_271 (N1206, N1010_t1, N938);
not NOT1_272 (N1207, N1013_t0);
nand NAND2_273 (N1208, N1013_t1, N942);
not NOT1_274 (N1209, N1016_t0);
nand NAND2_275 (N1210, N1016_t1, N946);
not NOT1_276 (N1211, N1019_t0);
nand NAND2_277 (N1212, N1019_t1, N950);
not NOT1_278 (N1213, N1022_t0);
nand NAND2_279 (N1214, N1022_t1, N954);
not NOT1_280 (N1215, N1025_t0);
nand NAND2_281 (N1216, N1025_t1, N958);
not NOT1_282 (N1217, N1028_t0);
not NOT1_283 (N1218, N959_t0);
not NOT1_284 (N1219, N1031_t0);
not NOT1_285 (N1220, N1034_t0);
nand NAND2_286 (N1221, N1034_t1, N968);
not NOT1_287 (N1222, N965_t0);
not NOT1_288 (N1223, N1037_t0);
nand NAND2_289 (N1224, N1037_t1, N972);
not NOT1_290 (N1225, N1040_t0);
nand NAND2_291 (N1226, N1040_t1, N976);
not NOT1_292 (N1227, N973_t0);
not NOT1_293 (N1228, N1043_t0);
nand NAND2_294 (N1229, N1043_t1, N980);
not NOT1_295 (N1230, N981_t0);
nand NAND2_296 (N1231, N981_t1, N984);
nand NAND2_297 (N1232, N1119, N1120);
nand NAND2_298 (N1235, N1121, N1122);
not NOT1_299 (N1238, N1046_t0);
nand NAND2_300 (N1239, N1046_t1, N997);
not NOT1_301 (N1240, N994_t0);
not NOT1_302 (N1241, N1049_t0);
nand NAND2_303 (N1242, N1049_t1, N1001);
nand NAND2_304 (N1243, N1128, N1129);
nand NAND2_305 (N1246, N1130, N1131);
nand NAND2_306 (N1249, N1132, N1133);
buf BUFF1_307 (N1252, N907_t0);
buf BUFF1_308 (N1255, N907_t1);
buf BUFF1_309 (N1258, N910_t0);
buf BUFF1_310 (N1261, N910_t1);
not NOT1_311 (N1264, N1150);
nand NAND2_312 (N1267, N631_t1, N1159);
nand NAND2_313 (N1309, N688_t1, N1205);
nand NAND2_314 (N1310, N691_t1, N1207);
nand NAND2_315 (N1311, N694_t1, N1209);
nand NAND2_316 (N1312, N697_t1, N1211);
nand NAND2_317 (N1313, N700_t1, N1213);
nand NAND2_318 (N1314, N703_t1, N1215);
nand NAND2_319 (N1315, N706_t1, N1220);
nand NAND2_320 (N1316, N709_t1, N1223);
nand NAND2_321 (N1317, N712_t1, N1225);
nand NAND2_322 (N1318, N715_t1, N1228);
not NOT1_323 (N1319, N1158);
nand NAND2_324 (N1322, N628_t1, N1230);
nand NAND2_325 (N1327, N730_t1, N1238);
nand NAND2_326 (N1328, N733_t1, N1241);
not NOT1_327 (N1334, N1162);
nand NAND2_328 (N1344, N1267, N1160);
nand NAND2_329 (N1345, N1249_t0, N894);
not NOT1_330 (N1346, N1249_t1);
not NOT1_331 (N1348, N1255_t0);
not NOT1_332 (N1349, N1252_t0);
not NOT1_333 (N1350, N1261_t0);
not NOT1_334 (N1351, N1258_t0);
nand NAND2_335 (N1352, N1309, N1206);
nand NAND2_336 (N1355, N1310, N1208);
nand NAND2_337 (N1358, N1311, N1210);
nand NAND2_338 (N1361, N1312, N1212);
nand NAND2_339 (N1364, N1313, N1214);
nand NAND2_340 (N1367, N1314, N1216);
nand NAND2_341 (N1370, N1315, N1221);
nand NAND2_342 (N1373, N1316, N1224);
nand NAND2_343 (N1376, N1317, N1226);
nand NAND2_344 (N1379, N1318, N1229);
nand NAND2_345 (N1383, N1322, N1231);
not NOT1_346 (N1386, N1232_t0);
nand NAND2_347 (N1387, N1232_t1, N990);
not NOT1_348 (N1388, N1235_t0);
nand NAND2_349 (N1389, N1235_t1, N993);
nand NAND2_350 (N1390, N1327, N1239);
nand NAND2_351 (N1393, N1328, N1242);
not NOT1_352 (N1396, N1243_t0);
nand NAND2_353 (N1397, N1243_t1, N1004);
not NOT1_354 (N1398, N1246_t0);
nand NAND2_355 (N1399, N1246_t1, N1007);
not NOT1_356 (N1409, N1319_t0);
nand NAND2_357 (N1412, N649_t1, N1346);
not NOT1_358 (N1413, N1334_t0);
buf BUFF1_359 (N1416, N1264_t0);
buf BUFF1_360 (N1419, N1264_t1);
nand NAND2_361 (N1433, N634_t1, N1386);
nand NAND2_362 (N1434, N637_t1, N1388);
nand NAND2_363 (N1438, N640_t1, N1396);
nand NAND2_364 (N1439, N646_t1, N1398);
not NOT1_365 (N1440, N1344);
nand NAND2_366 (N1443, N1355_t0, N1148);
not NOT1_367 (N1444, N1355_t1);
nand NAND2_368 (N1445, N1352_t0, N1149);
not NOT1_369 (N1446, N1352_t1);
nand NAND2_370 (N1447, N1358_t0, N1151);
not NOT1_371 (N1448, N1358_t1);
nand NAND2_372 (N1451, N1361_t0, N1152);
not NOT1_373 (N1452, N1361_t1);
nand NAND2_374 (N1453, N1367_t0, N1153);
not NOT1_375 (N1454, N1367_t1);
nand NAND2_376 (N1455, N1364_t0, N1154);
not NOT1_377 (N1456, N1364_t1);
nand NAND2_378 (N1457, N1373_t0, N1156);
not NOT1_379 (N1458, N1373_t1);
nand NAND2_380 (N1459, N1379_t0, N1157);
not NOT1_381 (N1460, N1379_t1);
not NOT1_382 (N1461, N1383_t0);
nand NAND2_383 (N1462, N1393_t0, N1161);
not NOT1_384 (N1463, N1393_t1);
nand NAND2_385 (N1464, N1345, N1412);
not NOT1_386 (N1468, N1370_t0);
nand NAND2_387 (N1469, N1370_t1, N1222);
not NOT1_388 (N1470, N1376_t0);
nand NAND2_389 (N1471, N1376_t1, N1227);
nand NAND2_390 (N1472, N1387, N1433);
not NOT1_391 (N1475, N1390_t0);
nand NAND2_392 (N1476, N1390_t1, N1240);
nand NAND2_393 (N1478, N1389, N1434);
nand NAND2_394 (N1481, N1399, N1439);
nand NAND2_395 (N1484, N1397, N1438);
nand NAND2_396 (N1487, N939_t1, N1444);
nand NAND2_397 (N1488, N935_t1, N1446);
nand NAND2_398 (N1489, N943_t1, N1448);
not NOT1_399 (N1490, N1419_t0);
not NOT1_400 (N1491, N1416_t0);
nand NAND2_401 (N1492, N947_t1, N1452);
nand NAND2_402 (N1493, N955_t1, N1454);
nand NAND2_403 (N1494, N951_t1, N1456);
nand NAND2_404 (N1495, N969_t1, N1458);
nand NAND2_405 (N1496, N977_t1, N1460);
nand NAND2_406 (N1498, N998_t1, N1463);
not NOT1_407 (N1499, N1440_t0);
nand NAND2_408 (N1500, N965_t1, N1468);
nand NAND2_409 (N1501, N973_t1, N1470);
nand NAND2_410 (N1504, N994_t1, N1475);
not NOT1_411 (N1510, N1464);
nand NAND2_412 (N1513, N1443, N1487);
nand NAND2_413 (N1514, N1445, N1488);
nand NAND2_414 (N1517, N1447, N1489);
nand NAND2_415 (N1520, N1451, N1492);
nand NAND2_416 (N1521, N1453, N1493);
nand NAND2_417 (N1522, N1455, N1494);
nand NAND2_418 (N1526, N1457, N1495);
nand NAND2_419 (N1527, N1459, N1496);
not NOT1_420 (N1528, N1472_t0);
nand NAND2_421 (N1529, N1462, N1498);
not NOT1_422 (N1530, N1478_t0);
not NOT1_423 (N1531, N1481_t0);
not NOT1_424 (N1532, N1484_t0);
nand NAND2_425 (N1534, N1471, N1501);
nand NAND2_426 (N1537, N1469, N1500);
nand NAND2_427 (N1540, N1476, N1504);
not NOT1_428 (N1546, N1513);
not NOT1_429 (N1554, N1521);
not NOT1_430 (N1557, N1526);
not NOT1_431 (N1561, N1520);
nand NAND2_432 (N1567, N1484_t1, N1531);
nand NAND2_433 (N1568, N1481_t1, N1532);
not NOT1_434 (N1569, N1510_t0);
not NOT1_435 (N1571, N1527);
not NOT1_436 (N1576, N1529);
buf BUFF1_437 (N1588, N1522_t0);
not NOT1_438 (N1591, N1534_t0);
not NOT1_439 (N1593, N1537_t0);
nand NAND2_440 (N1594, N1540_t0, N1530);
not NOT1_441 (N1595, N1540_t1);
nand NAND2_442 (N1596, N1567, N1568);
buf BUFF1_443 (N1600, N1517_t0);
buf BUFF1_444 (N1603, N1517_t1);
buf BUFF1_445 (N1606, N1522_t1);
buf BUFF1_446 (N1609, N1522_t2);
buf BUFF1_447 (N1612, N1514_t0);
buf BUFF1_448 (N1615, N1514_t1);
buf BUFF1_449 (N1620, N1557_t0);
buf BUFF1_450 (N1623, N1554_t0);
not NOT1_451 (N1635, N1571_t0);
nand NAND2_452 (N1636, N1478_t1, N1595);
nand NAND2_453 (N1638, N1576_t0, N1569);
not NOT1_454 (N1639, N1576_t1);
buf BUFF1_455 (N1640, N1561_t0);
buf BUFF1_456 (N1643, N1561_t1);
buf BUFF1_457 (N1647, N1546_t0);
buf BUFF1_458 (N1651, N1546_t1);
buf BUFF1_459 (N1658, N1554_t1);
buf BUFF1_460 (N1661, N1557_t1);
buf BUFF1_461 (N1664, N1557_t2);
nand NAND2_462 (N1671, N1596_t0, N893);
not NOT1_463 (N1672, N1596_t1);
not NOT1_464 (N1675, N1600_t0);
not NOT1_465 (N1677, N1603_t0);
nand NAND2_466 (N1678, N1606_t0, N1217);
not NOT1_467 (N1679, N1606_t1);
nand NAND2_468 (N1680, N1609_t0, N1219);
not NOT1_469 (N1681, N1609_t1);
not NOT1_470 (N1682, N1612_t0);
not NOT1_471 (N1683, N1615_t0);
nand NAND2_472 (N1685, N1594, N1636);
nand NAND2_473 (N1688, N1510_t1, N1639);
buf BUFF1_474 (N1697, N1588_t0);
buf BUFF1_475 (N1701, N1588_t1);
nand NAND2_476 (N1706, N643_t1, N1672);
not NOT1_477 (N1707, N1643_t0);
nand NAND2_478 (N1708, N1647_t0, N1675);
not NOT1_479 (N1709, N1647_t1);
nand NAND2_480 (N1710, N1651_t0, N1677);
not NOT1_481 (N1711, N1651_t1);
nand NAND2_482 (N1712, N1028_t1, N1679);
nand NAND2_483 (N1713, N1031_t1, N1681);
buf BUFF1_484 (N1714, N1620_t0);
buf BUFF1_485 (N1717, N1620_t1);
nand NAND2_486 (N1720, N1658_t0, N1593);
not NOT1_487 (N1721, N1658_t1);
nand NAND2_488 (N1723, N1638, N1688);
not NOT1_489 (N1727, N1661_t0);
not NOT1_490 (N1728, N1640_t0);
not NOT1_491 (N1730, N1664_t0);
buf BUFF1_492 (N1731, N1623_t0);
buf BUFF1_493 (N1734, N1623_t1);
nand NAND2_494 (N1740, N1685_t0, N1528);
not NOT1_495 (N1741, N1685_t1);
nand NAND2_496 (N1742, N1671, N1706);
nand NAND2_497 (N1746, N1600_t1, N1709);
nand NAND2_498 (N1747, N1603_t1, N1711);
nand NAND2_499 (N1748, N1678, N1712);
nand NAND2_500 (N1751, N1680, N1713);
nand NAND2_501 (N1759, N1537_t1, N1721);
not NOT1_502 (N1761, N1697_t0);
nand NAND2_503 (N1762, N1697_t1, N1727);
not NOT1_504 (N1763, N1701_t0);
nand NAND2_505 (N1764, N1701_t1, N1730);
not NOT1_506 (N1768, N1717_t0);
nand NAND2_507 (N1769, N1472_t1, N1741);
nand NAND2_508 (N1772, N1723_t0, N1413);
not NOT1_509 (N1773, N1723_t1);
nand NAND2_510 (N1774, N1708, N1746);
nand NAND2_511 (N1777, N1710, N1747);
not NOT1_512 (N1783, N1731_t0);
nand NAND2_513 (N1784, N1731_t1, N1682);
not NOT1_514 (N1785, N1714_t0);
not NOT1_515 (N1786, N1734_t0);
nand NAND2_516 (N1787, N1734_t1, N1683);
nand NAND2_517 (N1788, N1720, N1759);
nand NAND2_518 (N1791, N1661_t1, N1761);
nand NAND2_519 (N1792, N1664_t1, N1763);
nand NAND2_520 (N1795, N1751_t0, N1155);
not NOT1_521 (N1796, N1751_t1);
nand NAND2_522 (N1798, N1740, N1769);
nand NAND2_523 (N1801, N1334_t1, N1773);
nand NAND2_524 (N1802, N1742_t0, N290_t0);
not NOT1_525 (N1807, N1748_t0);
nand NAND2_526 (N1808, N1748_t1, N1218);
nand NAND2_527 (N1809, N1612_t1, N1783);
nand NAND2_528 (N1810, N1615_t1, N1786);
nand NAND2_529 (N1812, N1791, N1762);
nand NAND2_530 (N1815, N1792, N1764);
buf BUFF1_531 (N1818, N1742_t1);
nand NAND2_532 (N1821, N1777_t0, N1490);
not NOT1_533 (N1822, N1777_t1);
nand NAND2_534 (N1823, N1774_t0, N1491);
not NOT1_535 (N1824, N1774_t1);
nand NAND2_536 (N1825, N962_t1, N1796);
nand NAND2_537 (N1826, N1788_t0, N1409);
not NOT1_538 (N1827, N1788_t1);
nand NAND2_539 (N1830, N1772, N1801);
nand NAND2_540 (N1837, N959_t1, N1807);
nand NAND2_541 (N1838, N1809, N1784);
nand NAND2_542 (N1841, N1810, N1787);
nand NAND2_543 (N1848, N1419_t1, N1822);
nand NAND2_544 (N1849, N1416_t1, N1824);
nand NAND2_545 (N1850, N1795, N1825);
nand NAND2_546 (N1852, N1319_t1, N1827);
nand NAND2_547 (N1855, N1815_t0, N1707);
not NOT1_548 (N1856, N1815_t1);
not NOT1_549 (N1857, N1818_t0);
nand NAND2_550 (N1858, N1798_t0, N290_t1);
not NOT1_551 (N1864, N1812_t0);
nand NAND2_552 (N1865, N1812_t1, N1728);
buf BUFF1_553 (N1866, N1798_t1);
buf BUFF1_554 (N1869, N1802_t0);
buf BUFF1_555 (N1872, N1802_t1);
nand NAND2_556 (N1875, N1808, N1837);
nand NAND2_557 (N1878, N1821, N1848);
nand NAND2_558 (N1879, N1823, N1849);
nand NAND2_559 (N1882, N1841_t0, N1768);
not NOT1_560 (N1883, N1841_t1);
nand NAND2_561 (N1884, N1826, N1852);
nand NAND2_562 (N1885, N1643_t1, N1856);
nand NAND2_563 (N1889, N1830_t0, N290_t2);
not NOT1_564 (N1895, N1838_t0);
nand NAND2_565 (N1896, N1838_t1, N1785);
nand NAND2_566 (N1897, N1640_t1, N1864);
not NOT1_567 (N1898, N1850);
buf BUFF1_568 (N1902, N1830_t1);
not NOT1_569 (N1910, N1878);
nand NAND2_570 (N1911, N1717_t1, N1883);
not NOT1_571 (N1912, N1884);
nand NAND2_572 (N1913, N1855, N1885);
not NOT1_573 (N1915, N1866_t0);
nand NAND2_574 (N1919, N1872_t0, N919);
not NOT1_575 (N1920, N1872_t1);
nand NAND2_576 (N1921, N1869_t0, N920);
not NOT1_577 (N1922, N1869_t1);
not NOT1_578 (N1923, N1875_t0);
nand NAND2_579 (N1924, N1714_t1, N1895);
buf BUFF1_580 (N1927, N1858_t0);
buf BUFF1_581 (N1930, N1858_t1);
nand NAND2_582 (N1933, N1865, N1897);
nand NAND2_583 (N1936, N1882, N1911);
not NOT1_584 (N1937, N1898_t0);
not NOT1_585 (N1938, N1902_t0);
nand NAND2_586 (N1941, N679_t1, N1920);
nand NAND2_587 (N1942, N676_t1, N1922);
buf BUFF1_588 (N1944, N1879_t0);
not NOT1_589 (N1947, N1913);
buf BUFF1_590 (N1950, N1889_t0);
buf BUFF1_591 (N1953, N1889_t1);
buf BUFF1_592 (N1958, N1879_t1);
nand NAND2_593 (N1961, N1896, N1924);
and AND2_594 (N1965, N1910, N601);
and AND2_595 (N1968, N602, N1912);
nand NAND2_596 (N1975, N1930_t0, N917);
not NOT1_597 (N1976, N1930_t1);
nand NAND2_598 (N1977, N1927_t0, N918);
not NOT1_599 (N1978, N1927_t1);
nand NAND2_600 (N1979, N1919, N1941);
nand NAND2_601 (N1980, N1921, N1942);
not NOT1_602 (N1985, N1933_t0);
not NOT1_603 (N1987, N1936);
not NOT1_604 (N1999, N1944_t0);
nand NAND2_605 (N2000, N1944_t1, N1937);
not NOT1_606 (N2002, N1947_t0);
nand NAND2_607 (N2003, N1947_t1, N1499);
nand NAND2_608 (N2004, N1953_t0, N1350);
not NOT1_609 (N2005, N1953_t1);
nand NAND2_610 (N2006, N1950_t0, N1351);
not NOT1_611 (N2007, N1950_t1);
nand NAND2_612 (N2008, N673_t1, N1976);
nand NAND2_613 (N2009, N670_t1, N1978);
not NOT1_614 (N2012, N1979);
not NOT1_615 (N2013, N1958_t0);
nand NAND2_616 (N2014, N1958_t1, N1923);
not NOT1_617 (N2015, N1961_t0);
nand NAND2_618 (N2016, N1961_t1, N1635);
not NOT1_619 (N2018, N1965_t0);
not NOT1_620 (N2019, N1968_t0);
nand NAND2_621 (N2020, N1898_t1, N1999);
not NOT1_622 (N2021, N1987_t0);
nand NAND2_623 (N2022, N1987_t1, N1591);
nand NAND2_624 (N2023, N1440_t1, N2002);
nand NAND2_625 (N2024, N1261_t1, N2005);
nand NAND2_626 (N2025, N1258_t1, N2007);
nand NAND2_627 (N2026, N1975, N2008);
nand NAND2_628 (N2027, N1977, N2009);
not NOT1_629 (N2030, N1980_t0);
buf BUFF1_630 (N2033, N1980_t1);
nand NAND2_631 (N2036, N1875_t1, N2013);
nand NAND2_632 (N2037, N1571_t1, N2015);
nand NAND2_633 (N2038, N2020, N2000);
nand NAND2_634 (N2039, N1534_t1, N2021);
nand NAND2_635 (N2040, N2023, N2003);
nand NAND2_636 (N2041, N2004, N2024);
nand NAND2_637 (N2042, N2006, N2025);
not NOT1_638 (N2047, N2026);
nand NAND2_639 (N2052, N2036, N2014);
nand NAND2_640 (N2055, N2037, N2016);
not NOT1_641 (N2060, N2038);
nand NAND2_642 (N2061, N2039, N2022);
nand NAND2_643 (N2062, N2040, N290_t3);
not NOT1_644 (N2067, N2041);
not NOT1_645 (N2068, N2027_t0);
buf BUFF1_646 (N2071, N2027_t1);
not NOT1_647 (N2076, N2052_t0);
not NOT1_648 (N2077, N2055_t0);
nand NAND2_649 (N2078, N2060, N290_t4);
nand NAND2_650 (N2081, N2061, N290_t5);
not NOT1_651 (N2086, N2042_t0);
buf BUFF1_652 (N2089, N2042_t1);
and AND2_653 (N2104, N2030_t0, N2068_t0);
and AND2_654 (N2119, N2033_t0, N2068_t1);
and AND2_655 (N2129, N2030_t1, N2071_t0);
and AND2_656 (N2143, N2033_t1, N2071_t1);
buf BUFF1_657 (N2148, N2062_t0);
buf BUFF1_658 (N2151, N2062_t1);
buf BUFF1_659 (N2196, N2078_t0);
buf BUFF1_660 (N2199, N2078_t1);
buf BUFF1_661 (N2202, N2081_t0);
buf BUFF1_662 (N2205, N2081_t1);
nand NAND2_663 (N2214, N2151_t0, N915);
not NOT1_664 (N2215, N2151_t1);
nand NAND2_665 (N2216, N2148_t0, N916);
not NOT1_666 (N2217, N2148_t1);
nand NAND2_667 (N2222, N2199_t0, N1348);
not NOT1_668 (N2223, N2199_t1);
nand NAND2_669 (N2224, N2196_t0, N1349);
not NOT1_670 (N2225, N2196_t1);
nand NAND2_671 (N2226, N2205_t0, N913);
not NOT1_672 (N2227, N2205_t1);
nand NAND2_673 (N2228, N2202_t0, N914);
not NOT1_674 (N2229, N2202_t1);
nand NAND2_675 (N2230, N667_t1, N2215);
nand NAND2_676 (N2231, N664_t1, N2217);
nand NAND2_677 (N2232, N1255_t1, N2223);
nand NAND2_678 (N2233, N1252_t1, N2225);
nand NAND2_679 (N2234, N661_t1, N2227);
nand NAND2_680 (N2235, N658_t1, N2229);
nand NAND2_681 (N2236, N2214, N2230);
nand NAND2_682 (N2237, N2216, N2231);
nand NAND2_683 (N2240, N2222, N2232);
nand NAND2_684 (N2241, N2224, N2233);
nand NAND2_685 (N2244, N2226, N2234);
nand NAND2_686 (N2245, N2228, N2235);
not NOT1_687 (N2250, N2236);
not NOT1_688 (N2253, N2240);
not NOT1_689 (N2256, N2244);
not NOT1_690 (N2257, N2237_t0);
buf BUFF1_691 (N2260, N2237_t1);
not NOT1_692 (N2263, N2241_t0);
and AND2_693 (N2266, N1164_t0, N2241_t1);
not NOT1_694 (N2269, N2245_t0);
and AND2_695 (N2272, N1168_t0, N2245_t1);
nand NAND8_696 (N2279, N2067, N2012, N2047, N2250, N899_t2, N2256, N2253, N903_t2);
buf BUFF1_697 (N2286, N2266_t0);
buf BUFF1_698 (N2297, N2266_t1);
buf BUFF1_699 (N2315, N2272_t0);
buf BUFF1_700 (N2326, N2272_t1);
and AND2_701 (N2340, N2086_t0, N2257_t0);
and AND2_702 (N2353, N2089_t0, N2257_t1);
and AND2_703 (N2361, N2086_t1, N2260_t0);
and AND2_704 (N2375, N2089_t1, N2260_t1);
and AND4_705 (N2384, N338_t2, N2279_t0, N313_t0, N313);
and AND2_706 (N2385, N1163, N2263_t0);
and AND2_707 (N2386, N1164_t1, N2263_t1);
and AND2_708 (N2426, N1167, N2269_t0);
and AND2_709 (N2427, N1168_t1, N2269_t1);
nand NAND5_710 (N2537, N2286_t0, N2315_t0, N2361_t0, N2104_t0, N1171_t0);
nand NAND5_711 (N2540, N2286_t1, N2315_t1, N2340_t0, N2129_t0, N1171_t1);
nand NAND5_712 (N2543, N2286_t2, N2315_t2, N2340_t1, N2119_t0, N1171_t2);
nand NAND5_713 (N2546, N2286_t3, N2315_t3, N2353_t0, N2104_t1, N1171_t3);
nand NAND5_714 (N2549, N2297_t0, N2315_t4, N2375_t0, N2119_t1, N1188_t0);
nand NAND5_715 (N2552, N2297_t1, N2326_t0, N2361_t1, N2143_t0, N1188_t1);
nand NAND5_716 (N2555, N2297_t2, N2326_t1, N2375_t1, N2129_t1, N1188_t2);
and AND5_717 (N2558, N2286_t4, N2315_t5, N2361_t2, N2104_t2, N1171_t4);
and AND5_718 (N2561, N2286_t5, N2315_t6, N2340_t2, N2129_t2, N1171_t5);
and AND5_719 (N2564, N2286_t6, N2315_t7, N2340_t3, N2119_t2, N1171_t6);
and AND5_720 (N2567, N2286_t7, N2315_t8, N2353_t1, N2104_t3, N1171_t7);
and AND5_721 (N2570, N2297_t3, N2315_t9, N2375_t2, N2119_t3, N1188_t3);
and AND5_722 (N2573, N2297_t4, N2326_t2, N2361_t3, N2143_t1, N1188_t4);
and AND5_723 (N2576, N2297_t5, N2326_t3, N2375_t3, N2129_t3, N1188_t5);
nand NAND5_724 (N2594, N2286_t8, N2427_t0, N2361_t4, N2129_t4, N1171_t8);
nand NAND5_725 (N2597, N2297_t6, N2427_t1, N2361_t5, N2119_t4, N1171_t9);
nand NAND5_726 (N2600, N2297_t7, N2427_t2, N2375_t4, N2104_t4, N1171_t10);
nand NAND5_727 (N2603, N2297_t8, N2427_t3, N2340_t4, N2143_t2, N1171_t11);
nand NAND5_728 (N2606, N2297_t9, N2427_t4, N2353_t2, N2129_t5, N1188_t6);
nand NAND5_729 (N2611, N2386_t0, N2326_t4, N2361_t6, N2129_t6, N1188_t7);
nand NAND5_730 (N2614, N2386_t1, N2326_t5, N2361_t7, N2119_t5, N1188_t8);
nand NAND5_731 (N2617, N2386_t2, N2326_t6, N2375_t5, N2104_t5, N1188_t9);
nand NAND5_732 (N2620, N2386_t3, N2326_t7, N2353_t3, N2129_t7, N1188_t10);
nand NAND5_733 (N2627, N2297_t10, N2427_t5, N2340_t5, N2104_t6, N926_t0);
nand NAND5_734 (N2628, N2386_t4, N2326_t8, N2340_t6, N2104_t7, N926_t1);
nand NAND5_735 (N2629, N2386_t5, N2427_t6, N2361_t8, N2104_t8, N926_t2);
nand NAND5_736 (N2630, N2386_t6, N2427_t7, N2340_t7, N2129_t8, N926_t3);
nand NAND5_737 (N2631, N2386_t7, N2427_t8, N2340_t8, N2119_t6, N926_t4);
nand NAND5_738 (N2632, N2386_t8, N2427_t9, N2353_t4, N2104_t9, N926_t5);
nand NAND5_739 (N2633, N2386_t9, N2426, N2340_t9, N2104_t10, N926_t6);
nand NAND5_740 (N2634, N2385, N2427_t10, N2340_t10, N2104_t11, N926_t7);
and AND5_741 (N2639, N2286_t9, N2427_t11, N2361_t9, N2129_t9, N1171_t12);
and AND5_742 (N2642, N2297_t11, N2427_t12, N2361_t10, N2119_t7, N1171_t13);
and AND5_743 (N2645, N2297_t12, N2427_t13, N2375_t6, N2104_t12, N1171_t14);
and AND5_744 (N2648, N2297_t13, N2427_t14, N2340_t11, N2143_t3, N1171_t15);
and AND5_745 (N2651, N2297_t14, N2427_t15, N2353_t5, N2129_t10, N1188_t11);
and AND5_746 (N2655, N2386_t10, N2326_t9, N2361_t11, N2129_t11, N1188_t12);
and AND5_747 (N2658, N2386_t11, N2326_t10, N2361_t12, N2119_t8, N1188_t13);
and AND5_748 (N2661, N2386_t12, N2326_t11, N2375_t7, N2104_t13, N1188_t14);
and AND5_749 (N2664, N2386_t13, N2326_t12, N2353_t6, N2129_t12, N1188_t15);
nand NAND2_750 (N2669, N2558_t0, N534);
not NOT1_751 (N2670, N2558_t1);
nand NAND2_752 (N2671, N2561_t0, N535);
not NOT1_753 (N2672, N2561_t1);
nand NAND2_754 (N2673, N2564_t0, N536);
not NOT1_755 (N2674, N2564_t1);
nand NAND2_756 (N2675, N2567_t0, N537);
not NOT1_757 (N2676, N2567_t1);
nand NAND2_758 (N2682, N2570_t0, N543);
not NOT1_759 (N2683, N2570_t1);
nand NAND2_760 (N2688, N2573_t0, N548);
not NOT1_761 (N2689, N2573_t1);
nand NAND2_762 (N2690, N2576_t0, N549);
not NOT1_763 (N2691, N2576_t1);
and AND8_764 (N2710, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634);
nand NAND2_765 (N2720, N343_t1, N2670);
nand NAND2_766 (N2721, N346_t1, N2672);
nand NAND2_767 (N2722, N349_t1, N2674);
nand NAND2_768 (N2723, N352_t1, N2676);
nand NAND2_769 (N2724, N2639_t0, N538);
not NOT1_770 (N2725, N2639_t1);
nand NAND2_771 (N2726, N2642_t0, N539);
not NOT1_772 (N2727, N2642_t1);
nand NAND2_773 (N2728, N2645_t0, N540);
not NOT1_774 (N2729, N2645_t1);
nand NAND2_775 (N2730, N2648_t0, N541);
not NOT1_776 (N2731, N2648_t1);
nand NAND2_777 (N2732, N2651_t0, N542);
not NOT1_778 (N2733, N2651_t1);
nand NAND2_779 (N2734, N370_t1, N2683);
nand NAND2_780 (N2735, N2655_t0, N544);
not NOT1_781 (N2736, N2655_t1);
nand NAND2_782 (N2737, N2658_t0, N545);
not NOT1_783 (N2738, N2658_t1);
nand NAND2_784 (N2739, N2661_t0, N546);
not NOT1_785 (N2740, N2661_t1);
nand NAND2_786 (N2741, N2664_t0, N547);
not NOT1_787 (N2742, N2664_t1);
nand NAND2_788 (N2743, N385_t1, N2689);
nand NAND2_789 (N2744, N388_t1, N2691);
nand NAND8_790 (N2745, N2537_t0, N2540_t0, N2543_t0, N2546_t0, N2594_t0, N2597_t0, N2600_t0, N2603_t0);
nand NAND8_791 (N2746, N2606_t0, N2549_t0, N2611_t0, N2614_t0, N2617_t0, N2620_t0, N2552_t0, N2555_t0);
and AND8_792 (N2747, N2537_t1, N2540_t1, N2543_t1, N2546_t1, N2594_t1, N2597_t1, N2600_t1, N2603_t1);
and AND8_793 (N2750, N2606_t1, N2549_t1, N2611_t1, N2614_t1, N2617_t1, N2620_t1, N2552_t1, N2555_t1);
nand NAND2_794 (N2753, N2669, N2720);
nand NAND2_795 (N2754, N2671, N2721);
nand NAND2_796 (N2755, N2673, N2722);
nand NAND2_797 (N2756, N2675, N2723);
nand NAND2_798 (N2757, N355_t1, N2725);
nand NAND2_799 (N2758, N358_t1, N2727);
nand NAND2_800 (N2759, N361_t1, N2729);
nand NAND2_801 (N2760, N364_t1, N2731);
nand NAND2_802 (N2761, N367_t1, N2733);
nand NAND2_803 (N2762, N2682, N2734);
nand NAND2_804 (N2763, N373_t1, N2736);
nand NAND2_805 (N2764, N376_t1, N2738);
nand NAND2_806 (N2765, N379_t1, N2740);
nand NAND2_807 (N2766, N382_t1, N2742);
nand NAND2_808 (N2767, N2688, N2743);
nand NAND2_809 (N2768, N2690, N2744);
and AND2_810 (N2773, N2745, N275);
and AND2_811 (N2776, N2746, N276);
nand NAND2_812 (N2779, N2724, N2757);
nand NAND2_813 (N2780, N2726, N2758);
nand NAND2_814 (N2781, N2728, N2759);
nand NAND2_815 (N2782, N2730, N2760);
nand NAND2_816 (N2783, N2732, N2761);
nand NAND2_817 (N2784, N2735, N2763);
nand NAND2_818 (N2785, N2737, N2764);
nand NAND2_819 (N2786, N2739, N2765);
nand NAND2_820 (N2787, N2741, N2766);
and AND3_821 (N2788, N2747_t0, N2750_t0, N2710);
nand NAND2_822 (N2789, N2747_t1, N2750_t1);
and AND4_823 (N2800, N338_t3, N2279_t1, N99_t3, N2788);
nand NAND2_824 (N2807, N2773_t0, N2018);
not NOT1_825 (N2808, N2773_t1);
nand NAND2_826 (N2809, N2776_t0, N2019);
not NOT1_827 (N2810, N2776_t1);
nor NOR2_828 (N2811, N2384, N2800);
and AND3_829 (N2812, N897, N283_t0, N2789_t0);
and AND3_830 (N2815, N76_t1, N283_t1, N2789_t1);
and AND3_831 (N2818, N82_t1, N283_t2, N2789_t2);
and AND3_832 (N2821, N85_t1, N283_t3, N2789_t3);
and AND3_833 (N2824, N898, N283_t4, N2789_t4);
nand NAND2_834 (N2827, N1965_t1, N2808);
nand NAND2_835 (N2828, N1968_t1, N2810);
and AND3_836 (N2829, N79_t1, N283_t5, N2789_t5);
nand NAND2_837 (N2843, N2807, N2827);
nand NAND2_838 (N2846, N2809, N2828);
nand NAND2_839 (N2850, N2812_t0, N2076);
nand NAND2_840 (N2851, N2815_t0, N2077);
nand NAND2_841 (N2852, N2818_t0, N1915);
nand NAND2_842 (N2853, N2821_t0, N1857);
nand NAND2_843 (N2854, N2824_t0, N1938);
not NOT1_844 (N2857, N2812_t1);
not NOT1_845 (N2858, N2815_t1);
not NOT1_846 (N2859, N2818_t1);
not NOT1_847 (N2860, N2821_t1);
not NOT1_848 (N2861, N2824_t1);
not NOT1_849 (N2862, N2829_t0);
nand NAND2_850 (N2863, N2829_t1, N1985);
nand NAND2_851 (N2866, N2052_t1, N2857);
nand NAND2_852 (N2867, N2055_t1, N2858);
nand NAND2_853 (N2868, N1866_t1, N2859);
nand NAND2_854 (N2869, N1818_t1, N2860);
nand NAND2_855 (N2870, N1902_t1, N2861);
nand NAND2_856 (N2871, N2843_t0, N886);
not NOT1_857 (N2872, N2843_t1);
nand NAND2_858 (N2873, N2846_t0, N887);
not NOT1_859 (N2874, N2846_t1);
nand NAND2_860 (N2875, N1933_t1, N2862);
nand NAND2_861 (N2876, N2866, N2850);
nand NAND2_862 (N2877, N2867, N2851);
nand NAND2_863 (N2878, N2868, N2852);
nand NAND2_864 (N2879, N2869, N2853);
nand NAND2_865 (N2880, N2870, N2854);
nand NAND2_866 (N2881, N682_t1, N2872);
nand NAND2_867 (N2882, N685_t1, N2874);
nand NAND2_868 (N2883, N2875, N2863);
and AND2_869 (N2886, N2876, N550);
and AND2_870 (N2887, N551, N2877);
and AND2_871 (N2888, N553, N2878);
and AND2_872 (N2889, N2879, N554);
and AND2_873 (N2890, N555, N2880);
nand NAND2_874 (N2891, N2871, N2881);
nand NAND2_875 (N2892, N2873, N2882);
nand NAND2_876 (N2895, N2883_t0, N1461);
not NOT1_877 (N2896, N2883_t1);
nand NAND2_878 (N2897, N1383_t1, N2896);
nand NAND2_879 (N2898, N2895, N2897);
and AND2_880 (N2899, N2898, N552);

endmodule
