// Verilog
// c2670
// Ninputs 233
// Noutputs 140
// NtotalGates 1269
// BUFF1 272
// AND2 203
// NOT1 321
// AND4 11
// AND3 112
// NAND2 254
// OR2 51
// OR4 22
// NOR2 12
// AND5 7
// OR3 2
// OR5 2

module c2670f (INC,END,clk,rst,N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
              N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
              N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
              N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
              N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
              N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
              N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
              N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
              N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
              N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
              N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
              N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
              N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
              N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
              N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
              N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
              N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
              N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
              N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
              N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
              N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
              N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
              N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
              N216_I,N217_I,N218_I,N398,N400,N401,N419,N420,N456,N457,
              N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,
              N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,
              N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,
              N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,
              N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,
              N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,
              N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,
              N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,
              N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,
              N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,
              N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,
              N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,
              N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,
              N216_O,N217_O,N218_O);

input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
      N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
      N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
      N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
      N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
      N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
      N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
      N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
      N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
      N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
      N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
      N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
      N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
      N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
      N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
      N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
      N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
      N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
      N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
      N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
      N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
      N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
      N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
      N216_I,N217_I,N218_I;

output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,
       N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,
       N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,
       N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,
       N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,
       N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,
       N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,
       N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,
       N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,
       N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,
       N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,
       N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,
       N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,
       N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;

wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,
     N506,N509,N521,N533,N537,N543,N544,N547,N550,N562,
     N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,
     N612,N613,N625,N637,N643,N650,N651,N655,N659,N663,
     N667,N671,N675,N679,N683,N687,N693,N699,N705,N711,
     N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,
     N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,
     N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,
     N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,
     N1053,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1075,N1086,
     N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,
     N1127,N1128,N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,
     N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,N1173,N1178,
     N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,
     N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1219,N1222,N1225,
     N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,
     N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,
     N1353,N1354,N1355,N1395,N1396,N1397,N1398,N1399,N1422,N1423,
     N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,
     N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
     N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
     N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,
     N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,
     N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,
     N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
     N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
     N1549,N1550,N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,
     N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
     N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,
     N1612,N1615,N1619,N1624,N1628,N1631,N1634,N1637,N1642,N1647,
     N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,
     N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,
     N1808,N1809,N1810,N1811,N1813,N1814,N1815,N1822,N1823,N1824,
     N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,
     N1863,N1870,N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,
     N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
     N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,
     N1939,N1940,N1941,N1942,N1945,N1948,N1951,N1954,N1957,N1960,
     N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,
     N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,
     N2067,N2070,N2073,N2076,N2079,N2095,N2098,N2101,N2104,N2107,
     N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,
     N2144,N2147,N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,
     N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,N2188,N2191,
     N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,
     N2234,N2235,N2236,N2237,N2250,N2266,N2269,N2291,N2294,N2297,
     N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
     N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
     N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
     N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
     N2339,N2340,N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,
     N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,N2377,N2382,
     N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,
     N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2421,N2425,N2428,
     N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,
     N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,
     N2475,N2478,N2481,N2484,N2487,N2490,N2493,N2503,N2504,N2510,
     N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,
     N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,
     N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,N2610,N2611,
     N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,
     N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2638,N2645,N2646,
     N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,
     N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
     N2679,N2680,N2681,N2684,N2687,N2690,N2693,N2694,N2695,N2696,
     N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,
     N2709,N2710,N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,
     N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,N2773,N2774,
     N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,
     N2791,N2792,N2793,N2796,N2800,N2803,N2806,N2809,N2810,N2811,
     N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,
     N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,
     N2882,N2885,N2888,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
     N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,
     N2938,N2939,N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,
     N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,N3009,N3010,
     N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,
     N3037,N3039,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3053,
     N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,
     N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
     N3076,N3088,N3091,N3110,N3113,N3137,N3140,N3143,N3146,N3149,
     N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,
     N3178,N3180,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,
     N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,N3219,N3220,
     N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,
     N3256,N3259,N3262,N3265,N3268,N3271,N3274,N3277,N3281,N3282,
     N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,
     N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,
     N3321,N3324,N3327,N3330,N3333,N3334,N3335,N3336,N3337,N3340,
     N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,
     N3382,N3386,N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,
     N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,N3420,N3422,
     N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,
     N3459,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
     N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,
     N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
     N3509,N3510,N3511,N3512,N3513,N3515,N3517,N3522,N3525,N3528,
     N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,
     N3556,N3557,N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,
     N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,N3594,N3595,
     N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,
     N3622,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3640,N3644,
     N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,
     N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,
     N3720,N3721,N3722,N3723,N3726,N3727,N3728,N3729,N3730,N3731,
     N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,
     N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,N3780,N3790,
     N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,
     N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,
     N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,
     N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N1_t,N2_t,N3_t,N4_t,N5_t,N6_t,N7_t,N14_t,N15_t,N19_t,
     N20_t,N21_t,N22_t,N23_t,N24_t,N25_t,N26_t,N27_t,N28_t,N32_t,
     N33_t,N34_t,N35_t,N36_t,N43_t,N47_t,N48_t,N49_t,N50_t,N51_t,
     N52_t,N53_t,N54_t,N55_t,N56_t,N60_t,N61_t,N62_t,N63_t,N64_t,
     N65_t,N66_t,N67_t,N68_t,N72_t,N73_t,N74_t,N75_t,N76_t,N77_t,
     N78_t,N79_t,N80_t,N81_t,N85_t,N86_t,N87_t,N88_t,N89_t,N90_t,
     N91_t,N92_t,N93_t,N94_t,N95_t,N99_t,N100_t,N101_t,N102_t,N103_t,
     N104_t,N105_t,N106_t,N107_t,N111_t,N112_t,N113_t,N114_t,N115_t,N116_t,
     N117_t,N118_t,N119_t,N123_t,N124_t,N125_t,N126_t,N127_t,N128_t,N129_t,
     N130_t,N131_t,N135_t,N136_t,N137_t,N138_t,N139_t,N140_t,N141_t,N142_t,
     N230_t,N262_t,N143_I_t,N144_I_t,N145_I_t,N146_I_t,N147_I_t,N148_I_t,N149_I_t,N150_I_t,
     N151_I_t,N152_I_t,N153_I_t,N154_I_t,N155_I_t,N156_I_t,N157_I_t,N158_I_t,N159_I_t,N160_I_t,
     N161_I_t,N162_I_t,N163_I_t,N164_I_t,N165_I_t,N166_I_t,N167_I_t,N168_I_t,N169_I_t,N170_I_t,
     N171_I_t,N172_I_t,N173_I_t,N174_I_t,N175_I_t,N176_I_t,N177_I_t,N178_I_t,N179_I_t,N180_I_t,
     N181_I_t,N182_I_t,N183_I_t,N184_I_t,N185_I_t,N186_I_t,N187_I_t,N188_I_t,N189_I_t,N190_I_t,
     N191_I_t,N192_I_t,N193_I_t,N194_I_t,N195_I_t,N196_I_t,N197_I_t,N198_I_t,N199_I_t,N200_I_t,
     N201_I_t,N202_I_t,N203_I_t,N204_I_t,N205_I_t,N206_I_t,N207_I_t,N208_I_t,N209_I_t,N210_I_t,
     N211_I_t,N212_I_t,N213_I_t,N214_I_t,N215_I_t,N216_I_t,N217_I_t,N218_I_t;
wire N219_t0,N219_t1,N219_t2,N219_t3,N253_t0,N253_t1,N290_t0,N290_t1,N290_t2,
     N309_t0,N309_t1,N309_t2,N305_t0,N305_t1,N305_t2,N301_t0,N301_t1,N301_t2,N297_t0,
     N297_t1,N297_t2,N44_t0,N44_t1,N132_t0,N132_t1,N82_t0,N82_t1,N96_t0,N96_t1,
     N69_t0,N69_t1,N120_t0,N120_t1,N57_t0,N57_t1,N108_t0,N108_t1,N237_t0,N237_t1,
     N237_t2,N37_t0,N37_t1,N8_t0,N8_t1,N227_t0,N227_t1,N234_t0,N234_t1,N241_t0,
     N241_t1,N241_t2,N241_t3,N246_t0,N246_t1,N246_t2,N246_t3,N246_t4,N246_t5,N11_t0,
     N11_t1,N256_t0,N256_t1,N259_t0,N259_t1,N319_t0,N319_t1,N322_t0,N322_t1,N328_t0,
     N328_t1,N331_t0,N331_t1,N334_t0,N334_t1,N337_t0,N337_t1,N340_t0,N340_t1,N343_t0,
     N343_t1,N352_t0,N352_t1,N16_t0,N16_t1,N355_t0,N355_t1,N263_t0,N263_t1,N266_t0,
     N266_t1,N269_t0,N269_t1,N272_t0,N272_t1,N275_t0,N275_t1,N278_t0,N278_t1,N281_t0,
     N281_t1,N284_t0,N284_t1,N287_t0,N287_t1,N29_t0,N29_t1,N294_t0,N294_t1,N313_t0,
     N313_t1,N316_t0,N316_t1,N346_t0,N346_t1,N349_t0,N349_t1,N500_t0,N500_t1,N325_t0,
     N325_t1,N651_t0,N651_t1,N651_t2,N231_t0,N231_t1,N544_t0,N544_t1,N547_t0,N547_t1,
     N503_t0,N503_t1,N509_t0,N509_t1,N509_t2,N509_t3,N509_t4,N509_t5,N509_t6,N509_t7,
     N509_t8,N509_t9,N509_t10,N521_t0,N521_t1,N521_t2,N521_t3,N521_t4,N521_t5,N521_t6,
     N521_t7,N521_t8,N521_t9,N521_t10,N537_t0,N537_t1,N537_t2,N537_t3,N537_t4,N550_t0,
     N550_t1,N550_t2,N550_t3,N550_t4,N550_t5,N550_t6,N550_t7,N550_t8,N550_t9,N550_t10,
     N562_t0,N562_t1,N562_t2,N562_t3,N562_t4,N562_t5,N562_t6,N562_t7,N562_t8,N562_t9,
     N562_t10,N582_t0,N582_t1,N582_t2,N582_t3,N582_t4,N582_t5,N582_t6,N582_t7,N582_t8,
     N582_t9,N582_t10,N594_t0,N594_t1,N594_t2,N594_t3,N594_t4,N594_t5,N594_t6,N594_t7,
     N594_t8,N594_t9,N594_t10,N741_t0,N741_t1,N744_t0,N744_t1,N747_t0,N747_t1,N750_t0,
     N750_t1,N753_t0,N753_t1,N613_t0,N613_t1,N613_t2,N613_t3,N613_t4,N613_t5,N613_t6,
     N613_t7,N613_t8,N613_t9,N613_t10,N625_t0,N625_t1,N625_t2,N625_t3,N625_t4,N625_t5,
     N625_t6,N625_t7,N625_t8,N625_t9,N625_t10,N637_t0,N637_t1,N637_t2,N637_t3,N637_t4,
     N643_t0,N643_t1,N643_t2,N643_t3,N643_t4,N643_t5,N768_t0,N768_t1,N771_t0,N771_t1,
     N774_t0,N774_t1,N777_t0,N777_t1,N780_t0,N780_t1,N506_t0,N506_t1,N693_t0,N693_t1,
     N693_t2,N693_t3,N693_t4,N699_t0,N699_t1,N699_t2,N699_t3,N699_t4,N735_t0,N735_t1,
     N738_t0,N738_t1,N756_t0,N756_t1,N759_t0,N759_t1,N762_t0,N762_t1,N765_t0,N765_t1,
     N574_t0,N574_t1,N574_t2,N578_t0,N578_t1,N578_t2,N655_t0,N655_t1,N655_t2,N659_t0,
     N659_t1,N659_t2,N663_t0,N663_t1,N663_t2,N667_t0,N667_t1,N667_t2,N671_t0,N671_t1,
     N671_t2,N675_t0,N675_t1,N675_t2,N679_t0,N679_t1,N679_t2,N683_t0,N683_t1,N683_t2,
     N783_t0,N783_t1,N786_t0,N786_t1,N687_t0,N687_t1,N687_t2,N687_t3,N687_t4,N705_t0,
     N705_t1,N705_t2,N705_t3,N705_t4,N711_t0,N711_t1,N711_t2,N715_t0,N715_t1,N715_t2,
     N719_t0,N719_t1,N719_t2,N723_t0,N723_t1,N723_t2,N1034_t0,N1034_t1,N1042_t0,N1042_t1,
     N1042_t2,N1042_t3,N1042_t4,N1042_t5,N1042_t6,N1042_t7,N1042_t8,N1042_t9,N1053_t0,N1053_t1,
     N1053_t2,N1053_t3,N1053_t4,N1053_t5,N1053_t6,N1053_t7,N1053_t8,N1053_t9,N1075_t0,N1075_t1,
     N1075_t2,N1075_t3,N1075_t4,N1075_t5,N1075_t6,N1075_t7,N1075_t8,N1075_t9,N1086_t0,N1086_t1,
     N1086_t2,N1086_t3,N1086_t4,N1086_t5,N1086_t6,N1086_t7,N1086_t8,N1086_t9,N1102_t0,N1102_t1,
     N1102_t2,N1102_t3,N1102_t4,N1102_t5,N1102_t6,N1102_t7,N1102_t8,N1102_t9,N1113_t0,N1113_t1,
     N1113_t2,N1113_t3,N1113_t4,N1113_t5,N1113_t6,N1113_t7,N1113_t8,N1113_t9,N1129_t0,N1129_t1,
     N1129_t2,N1133_t0,N1133_t1,N1133_t2,N1137_t0,N1137_t1,N1219_t0,N1219_t1,N1222_t0,N1222_t1,
     N1225_t0,N1225_t1,N1228_t0,N1228_t1,N1231_t0,N1231_t1,N1234_t0,N1234_t1,N1237_t0,N1237_t1,
     N1240_t0,N1240_t1,N1243_t0,N1243_t1,N1246_t0,N1246_t1,N1146_t0,N1146_t1,N1146_t2,N1146_t3,
     N1146_t4,N1146_t5,N1146_t6,N1146_t7,N1146_t8,N1146_t9,N1157_t0,N1157_t1,N1157_t2,N1157_t3,
     N1157_t4,N1157_t5,N1157_t6,N1157_t7,N1157_t8,N1157_t9,N1173_t0,N1173_t1,N1173_t2,N1173_t3,
     N1178_t0,N1178_t1,N1178_t2,N1178_t3,N1178_t4,N1200_t0,N1200_t1,N1200_t2,N1200_t3,N1205_t0,
     N1205_t1,N1205_t2,N1205_t3,N1251_t0,N1251_t1,N1254_t0,N1254_t1,N1257_t0,N1257_t1,N1260_t0,
     N1260_t1,N1263_t0,N1263_t1,N1266_t0,N1266_t1,N1216_t0,N1216_t1,N1591_t0,N1591_t1,N1591_t2,
     N1591_t3,N1502_t0,N1502_t1,N1502_t2,N1506_t0,N1506_t1,N1506_t2,N1513_t0,N1513_t1,N1516_t0,
     N1516_t1,N1510_t0,N1510_t1,N1499_t0,N1499_t1,N1496_t0,N1496_t1,N1553_t0,N1553_t1,N1553_t2,
     N1557_t0,N1557_t1,N1557_t2,N1561_t0,N1561_t1,N1588_t0,N1588_t1,N1578_t0,N1578_t1,N1582_t0,
     N1582_t1,N1585_t0,N1585_t1,N1596_t0,N1596_t1,N1596_t2,N1606_t0,N1606_t1,N1606_t2,N1606_t3,
     N1606_t4,N1600_t0,N1600_t1,N1600_t2,N1600_t3,N1600_t4,N1642_t0,N1642_t1,N1642_t2,N1642_t3,
     N1647_t0,N1647_t1,N1647_t2,N1637_t0,N1637_t1,N1637_t2,N1637_t3,N1624_t0,N1624_t1,N1624_t2,
     N1619_t0,N1619_t1,N1619_t2,N1619_t3,N1615_t0,N1615_t1,N1615_t2,N496_t0,N496_t1,N224_t0,
     N224_t1,N1612_t0,N1612_t1,N1628_t0,N1628_t1,N1631_t0,N1631_t1,N1634_t0,N1634_t1,N727_t0,
     N727_t1,N1651_t0,N1651_t1,N1651_t2,N1651_t3,N730_t0,N730_t1,N1656_t0,N1656_t1,N1656_t2,
     N1686_t0,N1686_t1,N1686_t2,N1708_t0,N1708_t1,N1676_t0,N1676_t1,N1676_t2,N1676_t3,N1681_t0,
     N1681_t1,N1681_t2,N1681_t3,N1690_t0,N1690_t1,N533_t0,N533_t1,N533_t2,N1848_t0,N1848_t1,
     N1848_t2,N1852_t0,N1852_t1,N1852_t2,N1856_t0,N1856_t1,N1856_t2,N1856_t3,N1856_t4,N1856_t5,
     N1863_t0,N1863_t1,N1863_t2,N1863_t3,N1863_t4,N1863_t5,N1870_t0,N1870_t1,N1870_t2,N1870_t3,
     N1875_t0,N1875_t1,N1875_t2,N1875_t3,N1880_t0,N1880_t1,N1880_t2,N1880_t3,N1778_t0,N1778_t1,
     N1781_t0,N1781_t1,N1773_t0,N1773_t1,N1770_t0,N1770_t1,N1801_t0,N1801_t1,N1804_t0,N1804_t1,
     N1798_t0,N1798_t1,N1795_t0,N1795_t1,N1897_t0,N1897_t1,N1894_t0,N1894_t1,N40_t0,N40_t1,
     N1827_t0,N1827_t1,N1824_t0,N1824_t1,N1885_t0,N1885_t1,N1888_t0,N1888_t1,N1942_t0,N1942_t1,
     N1945_t0,N1945_t1,N1948_t0,N1948_t1,N1951_t0,N1951_t1,N1954_t0,N1954_t1,N1836_t0,N1836_t1,
     N1836_t2,N1836_t3,N1833_t0,N1833_t1,N1841_t0,N1841_t1,N1841_t2,N1841_t3,N1841_t4,N1841_t5,
     N1936_t0,N1936_t1,N1957_t0,N1957_t1,N1960_t0,N1960_t1,N1963_t0,N1963_t1,N1966_t0,N1966_t1,
     N2046_t0,N2046_t1,N2049_t0,N2049_t1,N2052_t0,N2052_t1,N2055_t0,N2055_t1,N2058_t0,N2058_t1,
     N2061_t0,N2061_t1,N2064_t0,N2064_t1,N2067_t0,N2067_t1,N2070_t0,N2070_t1,N2073_t0,N2073_t1,
     N2076_t0,N2076_t1,N2079_t0,N2079_t1,N2095_t0,N2095_t1,N2098_t0,N2098_t1,N2101_t0,N2101_t1,
     N2104_t0,N2104_t1,N2107_t0,N2107_t1,N2110_t0,N2110_t1,N2120_t0,N2120_t1,N2120_t2,N2120_t3,
     N2113_t0,N2113_t1,N2113_t2,N2113_t3,N2113_t4,N2185_t0,N2185_t1,N2188_t0,N2188_t1,N2191_t0,
     N2191_t1,N2194_t0,N2194_t1,N2201_t0,N2201_t1,N2204_t0,N2204_t1,N2207_t0,N2207_t1,N2210_t0,
     N2210_t1,N2213_t0,N2213_t1,N2266_t0,N2266_t1,N2269_t0,N2269_t1,N2219_t0,N2219_t1,N2216_t0,
     N2216_t1,N2128_t0,N2128_t1,N2128_t2,N2128_t3,N2128_t4,N2128_t5,N2135_t0,N2135_t1,N2135_t2,
     N2135_t3,N2135_t4,N2144_t0,N2144_t1,N2141_t0,N2141_t1,N2150_t0,N2150_t1,N2147_t0,N2147_t1,
     N2197_t0,N2197_t1,N2291_t0,N2291_t1,N2294_t0,N2294_t1,N2250_t0,N2250_t1,N2359_t0,N2359_t1,
     N2377_t0,N2377_t1,N2377_t2,N2377_t3,N1891_t0,N1891_t1,N2382_t0,N2382_t1,N2382_t2,N2434_t0,
     N2434_t1,N2437_t0,N2437_t1,N2368_t0,N2368_t1,N2368_t2,N2454_t0,N2454_t1,N2472_t0,N2472_t1,
     N2391_t0,N2391_t1,N2391_t2,N2395_t0,N2395_t1,N2395_t2,N2395_t3,N2521_t0,N2521_t1,N2475_t0,
     N2475_t1,N2478_t0,N2478_t1,N2481_t0,N2481_t1,N2484_t0,N2484_t1,N2417_t0,N2417_t1,N2417_t2,
     N2421_t0,N2421_t1,N2421_t2,N2425_t0,N2425_t1,N2493_t0,N2493_t1,N2440_t0,N2440_t1,N2443_t0,
     N2443_t1,N2446_t0,N2446_t1,N2449_t0,N2449_t1,N2457_t0,N2457_t1,N2460_t0,N2460_t1,N2463_t0,
     N2463_t1,N2466_t0,N2466_t1,N2469_t0,N2469_t1,N2487_t0,N2487_t1,N2490_t0,N2490_t1,N2534_t0,
     N2534_t1,N2531_t0,N2531_t1,N2537_t0,N2537_t1,N2540_t0,N2540_t1,N2638_t0,N2638_t1,N2638_t2,
     N2638_t3,N2613_t0,N2613_t1,N2613_t2,N2624_t0,N2624_t1,N2624_t2,N2646_t0,N2646_t1,N2646_t2,
     N2646_t3,N2603_t0,N2603_t1,N2603_t2,N2659_t0,N2659_t1,N2659_t2,N2687_t0,N2687_t1,N2690_t0,
     N2690_t1,N2684_t0,N2684_t1,N2681_t0,N2681_t1,N2703_t0,N2703_t1,N2729_t0,N2729_t1,N2729_t2,
     N2729_t3,N1037_t0,N1037_t1,N1037_t2,N1037_t3,N1070_t0,N1070_t1,N1070_t2,N1070_t3,N2738_t0,
     N2738_t1,N2738_t2,N2738_t3,N2817_t0,N2817_t1,N2841_t0,N2841_t1,N2826_t0,N2826_t1,N2796_t0,
     N2796_t1,N2796_t2,N2800_t0,N2800_t1,N2806_t0,N2806_t1,N2820_t0,N2820_t1,N2820_t2,N2820_t3,
     N2820_t4,N2831_t0,N2831_t1,N2831_t2,N2831_t3,N2831_t4,N2931_t0,N2931_t1,N2888_t0,N2888_t1,
     N2844_t0,N2844_t1,N2844_t2,N2844_t3,N2844_t4,N2854_t0,N2854_t1,N2854_t2,N2854_t3,N2859_t0,
     N2859_t1,N2859_t2,N2859_t3,N2859_t4,N2869_t0,N2869_t1,N2869_t2,N2869_t3,N2874_t0,N2874_t1,
     N2877_t0,N2877_t1,N2882_t0,N2882_t1,N2885_t0,N2885_t1,N1190_t0,N1190_t1,N1190_t2,N1190_t3,
     N2761_t0,N2761_t1,N2761_t2,N2761_t3,N1195_t0,N1195_t1,N1195_t2,N1195_t3,N2766_t0,N2766_t1,
     N2766_t2,N2766_t3,N2995_t0,N2995_t1,N2998_t0,N2998_t1,N3001_t0,N3001_t1,N3004_t0,N3004_t1,
     N2992_t0,N2992_t1,N2793_t0,N2793_t1,N2803_t0,N2803_t1,N2621_t0,N2621_t1,N3076_t0,N3076_t1,
     N3030_t0,N3030_t1,N3030_t2,N3030_t3,N3039_t0,N3039_t1,N3039_t2,N3039_t3,N3050_t0,N3050_t1,
     N3061_t0,N3061_t1,N2981_t0,N2981_t1,N2978_t0,N2978_t1,N2975_t0,N2975_t1,N2972_t0,N2972_t1,
     N2989_t0,N2989_t1,N2986_t0,N2986_t1,N3025_t0,N3025_t1,N3022_t0,N3022_t1,N3019_t0,N3019_t1,
     N3016_t0,N3016_t1,N3013_t0,N3013_t1,N3010_t0,N3010_t1,N3180_t0,N3180_t1,N3152_t0,N3152_t1,
     N3149_t0,N3149_t1,N3146_t0,N3146_t1,N3143_t0,N3143_t1,N3140_t0,N3140_t1,N3137_t0,N3137_t1,
     N3172_t0,N3172_t1,N3169_t0,N3169_t1,N3166_t0,N3166_t1,N3163_t0,N3163_t1,N3160_t0,N3160_t1,
     N3157_t0,N3157_t1,N3091_t0,N3091_t1,N3088_t0,N3088_t1,N3113_t0,N3113_t1,N3110_t0,N3110_t1,
     N3238_t0,N3238_t1,N3241_t0,N3241_t1,N3244_t0,N3244_t1,N3247_t0,N3247_t1,N3250_t0,N3250_t1,
     N3253_t0,N3253_t1,N3256_t0,N3256_t1,N3259_t0,N3259_t1,N3262_t0,N3262_t1,N3265_t0,N3265_t1,
     N3268_t0,N3268_t1,N3271_t0,N3271_t1,N3274_t0,N3274_t1,N3277_t0,N3277_t1,N3318_t0,N3318_t1,
     N3315_t0,N3315_t1,N3340_t0,N3340_t1,N3344_t0,N3344_t1,N3348_t0,N3348_t1,N3352_t0,N3352_t1,
     N3356_t0,N3356_t1,N3360_t0,N3360_t1,N3364_t0,N3364_t1,N3367_t0,N3367_t1,N3321_t0,N3321_t1,
     N3327_t0,N3327_t1,N3324_t0,N3324_t1,N3370_t0,N3370_t1,N3374_t0,N3374_t1,N3378_t0,N3378_t1,
     N3382_t0,N3382_t1,N3386_t0,N3386_t1,N3390_t0,N3390_t1,N3394_t0,N3394_t1,N3397_t0,N3397_t1,
     N3330_t0,N3330_t1,N3453_t0,N3453_t1,N3450_t0,N3450_t1,N3459_t0,N3459_t1,N3456_t0,N3456_t1,
     N3522_t0,N3522_t1,N3525_t0,N3525_t1,N3528_t0,N3528_t1,N3531_t0,N3531_t1,N800_t0,N800_t1,
     N3534_t0,N3534_t1,N3537_t0,N3537_t1,N3540_t0,N3540_t1,N3543_t0,N3543_t1,N3600_t0,N3600_t1,
     N3576_t0,N3576_t1,N3579_t0,N3579_t1,N3585_t0,N3585_t1,N3588_t0,N3588_t1,N3608_t0,N3608_t1,
     N3608_t2,N3612_t0,N3612_t1,N3603_t0,N3603_t1,N3603_t2,N3603_t3,N3616_t0,N3616_t1,N3616_t2,
     N3616_t3,N3616_t4,N3622_t0,N3622_t1,N3622_t2,N3622_t3,N3640_t0,N3640_t1,N3640_t2,N3644_t0,
     N3644_t1,N3635_t0,N3635_t1,N3635_t2,N3635_t3,N3648_t0,N3648_t1,N3648_t2,N3648_t3,N3648_t4,
     N3654_t0,N3654_t1,N3654_t2,N3654_t3,N3723_t0,N3723_t1,N3737_t0,N3737_t1,N3780_t0,N3780_t1,
     N3762_t0,N3762_t1,N3754_t0,N3754_t1,N3754_t2,N3758_t0,N3758_t1,N3790_t0,N3790_t1,N3775_t0,
     N3775_t1,N3767_t0,N3767_t1,N3767_t2,N3771_t0,N3771_t1,N3823_t0,N3823_t1,N3827_t0,N3827_t1,
     N3843_t0,N3843_t1,N3843_t2,N3840_t0,N3840_t1,N3852_t0,N3852_t1,N3859_t0,N3859_t1,N3864_t0,
     N3864_t1,N3870_t0,N3870_t1,N3877_t0,N3877_t1;
reg [1421:0] FEN;
fim PI_N1( .fault(fault), .net(N1), .FEN(FEN[0]), .op(N1_t) );
fim PI_N2( .fault(fault), .net(N2), .FEN(FEN[1]), .op(N2_t) );
fim PI_N3( .fault(fault), .net(N3), .FEN(FEN[2]), .op(N3_t) );
fim PI_N4( .fault(fault), .net(N4), .FEN(FEN[3]), .op(N4_t) );
fim PI_N5( .fault(fault), .net(N5), .FEN(FEN[4]), .op(N5_t) );
fim PI_N6( .fault(fault), .net(N6), .FEN(FEN[5]), .op(N6_t) );
fim PI_N7( .fault(fault), .net(N7), .FEN(FEN[6]), .op(N7_t) );
fim PI_N14( .fault(fault), .net(N14), .FEN(FEN[7]), .op(N14_t) );
fim PI_N15( .fault(fault), .net(N15), .FEN(FEN[8]), .op(N15_t) );
fim PI_N19( .fault(fault), .net(N19), .FEN(FEN[9]), .op(N19_t) );
fim PI_N20( .fault(fault), .net(N20), .FEN(FEN[10]), .op(N20_t) );
fim PI_N21( .fault(fault), .net(N21), .FEN(FEN[11]), .op(N21_t) );
fim PI_N22( .fault(fault), .net(N22), .FEN(FEN[12]), .op(N22_t) );
fim PI_N23( .fault(fault), .net(N23), .FEN(FEN[13]), .op(N23_t) );
fim PI_N24( .fault(fault), .net(N24), .FEN(FEN[14]), .op(N24_t) );
fim PI_N25( .fault(fault), .net(N25), .FEN(FEN[15]), .op(N25_t) );
fim PI_N26( .fault(fault), .net(N26), .FEN(FEN[16]), .op(N26_t) );
fim PI_N27( .fault(fault), .net(N27), .FEN(FEN[17]), .op(N27_t) );
fim PI_N28( .fault(fault), .net(N28), .FEN(FEN[18]), .op(N28_t) );
fim PI_N32( .fault(fault), .net(N32), .FEN(FEN[19]), .op(N32_t) );
fim PI_N33( .fault(fault), .net(N33), .FEN(FEN[20]), .op(N33_t) );
fim PI_N34( .fault(fault), .net(N34), .FEN(FEN[21]), .op(N34_t) );
fim PI_N35( .fault(fault), .net(N35), .FEN(FEN[22]), .op(N35_t) );
fim PI_N36( .fault(fault), .net(N36), .FEN(FEN[23]), .op(N36_t) );
fim PI_N43( .fault(fault), .net(N43), .FEN(FEN[24]), .op(N43_t) );
fim PI_N47( .fault(fault), .net(N47), .FEN(FEN[25]), .op(N47_t) );
fim PI_N48( .fault(fault), .net(N48), .FEN(FEN[26]), .op(N48_t) );
fim PI_N49( .fault(fault), .net(N49), .FEN(FEN[27]), .op(N49_t) );
fim PI_N50( .fault(fault), .net(N50), .FEN(FEN[28]), .op(N50_t) );
fim PI_N51( .fault(fault), .net(N51), .FEN(FEN[29]), .op(N51_t) );
fim PI_N52( .fault(fault), .net(N52), .FEN(FEN[30]), .op(N52_t) );
fim PI_N53( .fault(fault), .net(N53), .FEN(FEN[31]), .op(N53_t) );
fim PI_N54( .fault(fault), .net(N54), .FEN(FEN[32]), .op(N54_t) );
fim PI_N55( .fault(fault), .net(N55), .FEN(FEN[33]), .op(N55_t) );
fim PI_N56( .fault(fault), .net(N56), .FEN(FEN[34]), .op(N56_t) );
fim PI_N60( .fault(fault), .net(N60), .FEN(FEN[35]), .op(N60_t) );
fim PI_N61( .fault(fault), .net(N61), .FEN(FEN[36]), .op(N61_t) );
fim PI_N62( .fault(fault), .net(N62), .FEN(FEN[37]), .op(N62_t) );
fim PI_N63( .fault(fault), .net(N63), .FEN(FEN[38]), .op(N63_t) );
fim PI_N64( .fault(fault), .net(N64), .FEN(FEN[39]), .op(N64_t) );
fim PI_N65( .fault(fault), .net(N65), .FEN(FEN[40]), .op(N65_t) );
fim PI_N66( .fault(fault), .net(N66), .FEN(FEN[41]), .op(N66_t) );
fim PI_N67( .fault(fault), .net(N67), .FEN(FEN[42]), .op(N67_t) );
fim PI_N68( .fault(fault), .net(N68), .FEN(FEN[43]), .op(N68_t) );
fim PI_N72( .fault(fault), .net(N72), .FEN(FEN[44]), .op(N72_t) );
fim PI_N73( .fault(fault), .net(N73), .FEN(FEN[45]), .op(N73_t) );
fim PI_N74( .fault(fault), .net(N74), .FEN(FEN[46]), .op(N74_t) );
fim PI_N75( .fault(fault), .net(N75), .FEN(FEN[47]), .op(N75_t) );
fim PI_N76( .fault(fault), .net(N76), .FEN(FEN[48]), .op(N76_t) );
fim PI_N77( .fault(fault), .net(N77), .FEN(FEN[49]), .op(N77_t) );
fim PI_N78( .fault(fault), .net(N78), .FEN(FEN[50]), .op(N78_t) );
fim PI_N79( .fault(fault), .net(N79), .FEN(FEN[51]), .op(N79_t) );
fim PI_N80( .fault(fault), .net(N80), .FEN(FEN[52]), .op(N80_t) );
fim PI_N81( .fault(fault), .net(N81), .FEN(FEN[53]), .op(N81_t) );
fim PI_N85( .fault(fault), .net(N85), .FEN(FEN[54]), .op(N85_t) );
fim PI_N86( .fault(fault), .net(N86), .FEN(FEN[55]), .op(N86_t) );
fim PI_N87( .fault(fault), .net(N87), .FEN(FEN[56]), .op(N87_t) );
fim PI_N88( .fault(fault), .net(N88), .FEN(FEN[57]), .op(N88_t) );
fim PI_N89( .fault(fault), .net(N89), .FEN(FEN[58]), .op(N89_t) );
fim PI_N90( .fault(fault), .net(N90), .FEN(FEN[59]), .op(N90_t) );
fim PI_N91( .fault(fault), .net(N91), .FEN(FEN[60]), .op(N91_t) );
fim PI_N92( .fault(fault), .net(N92), .FEN(FEN[61]), .op(N92_t) );
fim PI_N93( .fault(fault), .net(N93), .FEN(FEN[62]), .op(N93_t) );
fim PI_N94( .fault(fault), .net(N94), .FEN(FEN[63]), .op(N94_t) );
fim PI_N95( .fault(fault), .net(N95), .FEN(FEN[64]), .op(N95_t) );
fim PI_N99( .fault(fault), .net(N99), .FEN(FEN[65]), .op(N99_t) );
fim PI_N100( .fault(fault), .net(N100), .FEN(FEN[66]), .op(N100_t) );
fim PI_N101( .fault(fault), .net(N101), .FEN(FEN[67]), .op(N101_t) );
fim PI_N102( .fault(fault), .net(N102), .FEN(FEN[68]), .op(N102_t) );
fim PI_N103( .fault(fault), .net(N103), .FEN(FEN[69]), .op(N103_t) );
fim PI_N104( .fault(fault), .net(N104), .FEN(FEN[70]), .op(N104_t) );
fim PI_N105( .fault(fault), .net(N105), .FEN(FEN[71]), .op(N105_t) );
fim PI_N106( .fault(fault), .net(N106), .FEN(FEN[72]), .op(N106_t) );
fim PI_N107( .fault(fault), .net(N107), .FEN(FEN[73]), .op(N107_t) );
fim PI_N111( .fault(fault), .net(N111), .FEN(FEN[74]), .op(N111_t) );
fim PI_N112( .fault(fault), .net(N112), .FEN(FEN[75]), .op(N112_t) );
fim PI_N113( .fault(fault), .net(N113), .FEN(FEN[76]), .op(N113_t) );
fim PI_N114( .fault(fault), .net(N114), .FEN(FEN[77]), .op(N114_t) );
fim PI_N115( .fault(fault), .net(N115), .FEN(FEN[78]), .op(N115_t) );
fim PI_N116( .fault(fault), .net(N116), .FEN(FEN[79]), .op(N116_t) );
fim PI_N117( .fault(fault), .net(N117), .FEN(FEN[80]), .op(N117_t) );
fim PI_N118( .fault(fault), .net(N118), .FEN(FEN[81]), .op(N118_t) );
fim PI_N119( .fault(fault), .net(N119), .FEN(FEN[82]), .op(N119_t) );
fim PI_N123( .fault(fault), .net(N123), .FEN(FEN[83]), .op(N123_t) );
fim PI_N124( .fault(fault), .net(N124), .FEN(FEN[84]), .op(N124_t) );
fim PI_N125( .fault(fault), .net(N125), .FEN(FEN[85]), .op(N125_t) );
fim PI_N126( .fault(fault), .net(N126), .FEN(FEN[86]), .op(N126_t) );
fim PI_N127( .fault(fault), .net(N127), .FEN(FEN[87]), .op(N127_t) );
fim PI_N128( .fault(fault), .net(N128), .FEN(FEN[88]), .op(N128_t) );
fim PI_N129( .fault(fault), .net(N129), .FEN(FEN[89]), .op(N129_t) );
fim PI_N130( .fault(fault), .net(N130), .FEN(FEN[90]), .op(N130_t) );
fim PI_N131( .fault(fault), .net(N131), .FEN(FEN[91]), .op(N131_t) );
fim PI_N135( .fault(fault), .net(N135), .FEN(FEN[92]), .op(N135_t) );
fim PI_N136( .fault(fault), .net(N136), .FEN(FEN[93]), .op(N136_t) );
fim PI_N137( .fault(fault), .net(N137), .FEN(FEN[94]), .op(N137_t) );
fim PI_N138( .fault(fault), .net(N138), .FEN(FEN[95]), .op(N138_t) );
fim PI_N139( .fault(fault), .net(N139), .FEN(FEN[96]), .op(N139_t) );
fim PI_N140( .fault(fault), .net(N140), .FEN(FEN[97]), .op(N140_t) );
fim PI_N141( .fault(fault), .net(N141), .FEN(FEN[98]), .op(N141_t) );
fim PI_N142( .fault(fault), .net(N142), .FEN(FEN[99]), .op(N142_t) );
fim PI_N230( .fault(fault), .net(N230), .FEN(FEN[100]), .op(N230_t) );
fim PI_N262( .fault(fault), .net(N262), .FEN(FEN[101]), .op(N262_t) );
fim PI_N143_I( .fault(fault), .net(N143_I), .FEN(FEN[102]), .op(N143_I_t) );
fim PI_N144_I( .fault(fault), .net(N144_I), .FEN(FEN[103]), .op(N144_I_t) );
fim PI_N145_I( .fault(fault), .net(N145_I), .FEN(FEN[104]), .op(N145_I_t) );
fim PI_N146_I( .fault(fault), .net(N146_I), .FEN(FEN[105]), .op(N146_I_t) );
fim PI_N147_I( .fault(fault), .net(N147_I), .FEN(FEN[106]), .op(N147_I_t) );
fim PI_N148_I( .fault(fault), .net(N148_I), .FEN(FEN[107]), .op(N148_I_t) );
fim PI_N149_I( .fault(fault), .net(N149_I), .FEN(FEN[108]), .op(N149_I_t) );
fim PI_N150_I( .fault(fault), .net(N150_I), .FEN(FEN[109]), .op(N150_I_t) );
fim PI_N151_I( .fault(fault), .net(N151_I), .FEN(FEN[110]), .op(N151_I_t) );
fim PI_N152_I( .fault(fault), .net(N152_I), .FEN(FEN[111]), .op(N152_I_t) );
fim PI_N153_I( .fault(fault), .net(N153_I), .FEN(FEN[112]), .op(N153_I_t) );
fim PI_N154_I( .fault(fault), .net(N154_I), .FEN(FEN[113]), .op(N154_I_t) );
fim PI_N155_I( .fault(fault), .net(N155_I), .FEN(FEN[114]), .op(N155_I_t) );
fim PI_N156_I( .fault(fault), .net(N156_I), .FEN(FEN[115]), .op(N156_I_t) );
fim PI_N157_I( .fault(fault), .net(N157_I), .FEN(FEN[116]), .op(N157_I_t) );
fim PI_N158_I( .fault(fault), .net(N158_I), .FEN(FEN[117]), .op(N158_I_t) );
fim PI_N159_I( .fault(fault), .net(N159_I), .FEN(FEN[118]), .op(N159_I_t) );
fim PI_N160_I( .fault(fault), .net(N160_I), .FEN(FEN[119]), .op(N160_I_t) );
fim PI_N161_I( .fault(fault), .net(N161_I), .FEN(FEN[120]), .op(N161_I_t) );
fim PI_N162_I( .fault(fault), .net(N162_I), .FEN(FEN[121]), .op(N162_I_t) );
fim PI_N163_I( .fault(fault), .net(N163_I), .FEN(FEN[122]), .op(N163_I_t) );
fim PI_N164_I( .fault(fault), .net(N164_I), .FEN(FEN[123]), .op(N164_I_t) );
fim PI_N165_I( .fault(fault), .net(N165_I), .FEN(FEN[124]), .op(N165_I_t) );
fim PI_N166_I( .fault(fault), .net(N166_I), .FEN(FEN[125]), .op(N166_I_t) );
fim PI_N167_I( .fault(fault), .net(N167_I), .FEN(FEN[126]), .op(N167_I_t) );
fim PI_N168_I( .fault(fault), .net(N168_I), .FEN(FEN[127]), .op(N168_I_t) );
fim PI_N169_I( .fault(fault), .net(N169_I), .FEN(FEN[128]), .op(N169_I_t) );
fim PI_N170_I( .fault(fault), .net(N170_I), .FEN(FEN[129]), .op(N170_I_t) );
fim PI_N171_I( .fault(fault), .net(N171_I), .FEN(FEN[130]), .op(N171_I_t) );
fim PI_N172_I( .fault(fault), .net(N172_I), .FEN(FEN[131]), .op(N172_I_t) );
fim PI_N173_I( .fault(fault), .net(N173_I), .FEN(FEN[132]), .op(N173_I_t) );
fim PI_N174_I( .fault(fault), .net(N174_I), .FEN(FEN[133]), .op(N174_I_t) );
fim PI_N175_I( .fault(fault), .net(N175_I), .FEN(FEN[134]), .op(N175_I_t) );
fim PI_N176_I( .fault(fault), .net(N176_I), .FEN(FEN[135]), .op(N176_I_t) );
fim PI_N177_I( .fault(fault), .net(N177_I), .FEN(FEN[136]), .op(N177_I_t) );
fim PI_N178_I( .fault(fault), .net(N178_I), .FEN(FEN[137]), .op(N178_I_t) );
fim PI_N179_I( .fault(fault), .net(N179_I), .FEN(FEN[138]), .op(N179_I_t) );
fim PI_N180_I( .fault(fault), .net(N180_I), .FEN(FEN[139]), .op(N180_I_t) );
fim PI_N181_I( .fault(fault), .net(N181_I), .FEN(FEN[140]), .op(N181_I_t) );
fim PI_N182_I( .fault(fault), .net(N182_I), .FEN(FEN[141]), .op(N182_I_t) );
fim PI_N183_I( .fault(fault), .net(N183_I), .FEN(FEN[142]), .op(N183_I_t) );
fim PI_N184_I( .fault(fault), .net(N184_I), .FEN(FEN[143]), .op(N184_I_t) );
fim PI_N185_I( .fault(fault), .net(N185_I), .FEN(FEN[144]), .op(N185_I_t) );
fim PI_N186_I( .fault(fault), .net(N186_I), .FEN(FEN[145]), .op(N186_I_t) );
fim PI_N187_I( .fault(fault), .net(N187_I), .FEN(FEN[146]), .op(N187_I_t) );
fim PI_N188_I( .fault(fault), .net(N188_I), .FEN(FEN[147]), .op(N188_I_t) );
fim PI_N189_I( .fault(fault), .net(N189_I), .FEN(FEN[148]), .op(N189_I_t) );
fim PI_N190_I( .fault(fault), .net(N190_I), .FEN(FEN[149]), .op(N190_I_t) );
fim PI_N191_I( .fault(fault), .net(N191_I), .FEN(FEN[150]), .op(N191_I_t) );
fim PI_N192_I( .fault(fault), .net(N192_I), .FEN(FEN[151]), .op(N192_I_t) );
fim PI_N193_I( .fault(fault), .net(N193_I), .FEN(FEN[152]), .op(N193_I_t) );
fim PI_N194_I( .fault(fault), .net(N194_I), .FEN(FEN[153]), .op(N194_I_t) );
fim PI_N195_I( .fault(fault), .net(N195_I), .FEN(FEN[154]), .op(N195_I_t) );
fim PI_N196_I( .fault(fault), .net(N196_I), .FEN(FEN[155]), .op(N196_I_t) );
fim PI_N197_I( .fault(fault), .net(N197_I), .FEN(FEN[156]), .op(N197_I_t) );
fim PI_N198_I( .fault(fault), .net(N198_I), .FEN(FEN[157]), .op(N198_I_t) );
fim PI_N199_I( .fault(fault), .net(N199_I), .FEN(FEN[158]), .op(N199_I_t) );
fim PI_N200_I( .fault(fault), .net(N200_I), .FEN(FEN[159]), .op(N200_I_t) );
fim PI_N201_I( .fault(fault), .net(N201_I), .FEN(FEN[160]), .op(N201_I_t) );
fim PI_N202_I( .fault(fault), .net(N202_I), .FEN(FEN[161]), .op(N202_I_t) );
fim PI_N203_I( .fault(fault), .net(N203_I), .FEN(FEN[162]), .op(N203_I_t) );
fim PI_N204_I( .fault(fault), .net(N204_I), .FEN(FEN[163]), .op(N204_I_t) );
fim PI_N205_I( .fault(fault), .net(N205_I), .FEN(FEN[164]), .op(N205_I_t) );
fim PI_N206_I( .fault(fault), .net(N206_I), .FEN(FEN[165]), .op(N206_I_t) );
fim PI_N207_I( .fault(fault), .net(N207_I), .FEN(FEN[166]), .op(N207_I_t) );
fim PI_N208_I( .fault(fault), .net(N208_I), .FEN(FEN[167]), .op(N208_I_t) );
fim PI_N209_I( .fault(fault), .net(N209_I), .FEN(FEN[168]), .op(N209_I_t) );
fim PI_N210_I( .fault(fault), .net(N210_I), .FEN(FEN[169]), .op(N210_I_t) );
fim PI_N211_I( .fault(fault), .net(N211_I), .FEN(FEN[170]), .op(N211_I_t) );
fim PI_N212_I( .fault(fault), .net(N212_I), .FEN(FEN[171]), .op(N212_I_t) );
fim PI_N213_I( .fault(fault), .net(N213_I), .FEN(FEN[172]), .op(N213_I_t) );
fim PI_N214_I( .fault(fault), .net(N214_I), .FEN(FEN[173]), .op(N214_I_t) );
fim PI_N215_I( .fault(fault), .net(N215_I), .FEN(FEN[174]), .op(N215_I_t) );
fim PI_N216_I( .fault(fault), .net(N216_I), .FEN(FEN[175]), .op(N216_I_t) );
fim PI_N217_I( .fault(fault), .net(N217_I), .FEN(FEN[176]), .op(N217_I_t) );
fim PI_N218_I( .fault(fault), .net(N218_I), .FEN(FEN[177]), .op(N218_I_t) );
fim FAN_N219_0 ( .fault(fault), .net(N219), .FEN(FEN[178]), .op(N219_t0) );
fim FAN_N219_1 ( .fault(fault), .net(N219), .FEN(FEN[179]), .op(N219_t1) );
fim FAN_N219_2 ( .fault(fault), .net(N219), .FEN(FEN[180]), .op(N219_t2) );
fim FAN_N219_3 ( .fault(fault), .net(N219), .FEN(FEN[181]), .op(N219_t3) );
fim FAN_N253_0 ( .fault(fault), .net(N253), .FEN(FEN[182]), .op(N253_t0) );
fim FAN_N253_1 ( .fault(fault), .net(N253), .FEN(FEN[183]), .op(N253_t1) );
fim FAN_N290_0 ( .fault(fault), .net(N290), .FEN(FEN[184]), .op(N290_t0) );
fim FAN_N290_1 ( .fault(fault), .net(N290), .FEN(FEN[185]), .op(N290_t1) );
fim FAN_N290_2 ( .fault(fault), .net(N290), .FEN(FEN[186]), .op(N290_t2) );
fim FAN_N309_0 ( .fault(fault), .net(N309), .FEN(FEN[187]), .op(N309_t0) );
fim FAN_N309_1 ( .fault(fault), .net(N309), .FEN(FEN[188]), .op(N309_t1) );
fim FAN_N309_2 ( .fault(fault), .net(N309), .FEN(FEN[189]), .op(N309_t2) );
fim FAN_N305_0 ( .fault(fault), .net(N305), .FEN(FEN[190]), .op(N305_t0) );
fim FAN_N305_1 ( .fault(fault), .net(N305), .FEN(FEN[191]), .op(N305_t1) );
fim FAN_N305_2 ( .fault(fault), .net(N305), .FEN(FEN[192]), .op(N305_t2) );
fim FAN_N301_0 ( .fault(fault), .net(N301), .FEN(FEN[193]), .op(N301_t0) );
fim FAN_N301_1 ( .fault(fault), .net(N301), .FEN(FEN[194]), .op(N301_t1) );
fim FAN_N301_2 ( .fault(fault), .net(N301), .FEN(FEN[195]), .op(N301_t2) );
fim FAN_N297_0 ( .fault(fault), .net(N297), .FEN(FEN[196]), .op(N297_t0) );
fim FAN_N297_1 ( .fault(fault), .net(N297), .FEN(FEN[197]), .op(N297_t1) );
fim FAN_N297_2 ( .fault(fault), .net(N297), .FEN(FEN[198]), .op(N297_t2) );
fim FAN_N44_0 ( .fault(fault), .net(N44), .FEN(FEN[199]), .op(N44_t0) );
fim FAN_N44_1 ( .fault(fault), .net(N44), .FEN(FEN[200]), .op(N44_t1) );
fim FAN_N132_0 ( .fault(fault), .net(N132), .FEN(FEN[201]), .op(N132_t0) );
fim FAN_N132_1 ( .fault(fault), .net(N132), .FEN(FEN[202]), .op(N132_t1) );
fim FAN_N82_0 ( .fault(fault), .net(N82), .FEN(FEN[203]), .op(N82_t0) );
fim FAN_N82_1 ( .fault(fault), .net(N82), .FEN(FEN[204]), .op(N82_t1) );
fim FAN_N96_0 ( .fault(fault), .net(N96), .FEN(FEN[205]), .op(N96_t0) );
fim FAN_N96_1 ( .fault(fault), .net(N96), .FEN(FEN[206]), .op(N96_t1) );
fim FAN_N69_0 ( .fault(fault), .net(N69), .FEN(FEN[207]), .op(N69_t0) );
fim FAN_N69_1 ( .fault(fault), .net(N69), .FEN(FEN[208]), .op(N69_t1) );
fim FAN_N120_0 ( .fault(fault), .net(N120), .FEN(FEN[209]), .op(N120_t0) );
fim FAN_N120_1 ( .fault(fault), .net(N120), .FEN(FEN[210]), .op(N120_t1) );
fim FAN_N57_0 ( .fault(fault), .net(N57), .FEN(FEN[211]), .op(N57_t0) );
fim FAN_N57_1 ( .fault(fault), .net(N57), .FEN(FEN[212]), .op(N57_t1) );
fim FAN_N108_0 ( .fault(fault), .net(N108), .FEN(FEN[213]), .op(N108_t0) );
fim FAN_N108_1 ( .fault(fault), .net(N108), .FEN(FEN[214]), .op(N108_t1) );
fim FAN_N237_0 ( .fault(fault), .net(N237), .FEN(FEN[215]), .op(N237_t0) );
fim FAN_N237_1 ( .fault(fault), .net(N237), .FEN(FEN[216]), .op(N237_t1) );
fim FAN_N237_2 ( .fault(fault), .net(N237), .FEN(FEN[217]), .op(N237_t2) );
fim FAN_N37_0 ( .fault(fault), .net(N37), .FEN(FEN[218]), .op(N37_t0) );
fim FAN_N37_1 ( .fault(fault), .net(N37), .FEN(FEN[219]), .op(N37_t1) );
fim FAN_N8_0 ( .fault(fault), .net(N8), .FEN(FEN[220]), .op(N8_t0) );
fim FAN_N8_1 ( .fault(fault), .net(N8), .FEN(FEN[221]), .op(N8_t1) );
fim FAN_N227_0 ( .fault(fault), .net(N227), .FEN(FEN[222]), .op(N227_t0) );
fim FAN_N227_1 ( .fault(fault), .net(N227), .FEN(FEN[223]), .op(N227_t1) );
fim FAN_N234_0 ( .fault(fault), .net(N234), .FEN(FEN[224]), .op(N234_t0) );
fim FAN_N234_1 ( .fault(fault), .net(N234), .FEN(FEN[225]), .op(N234_t1) );
fim FAN_N241_0 ( .fault(fault), .net(N241), .FEN(FEN[226]), .op(N241_t0) );
fim FAN_N241_1 ( .fault(fault), .net(N241), .FEN(FEN[227]), .op(N241_t1) );
fim FAN_N241_2 ( .fault(fault), .net(N241), .FEN(FEN[228]), .op(N241_t2) );
fim FAN_N241_3 ( .fault(fault), .net(N241), .FEN(FEN[229]), .op(N241_t3) );
fim FAN_N246_0 ( .fault(fault), .net(N246), .FEN(FEN[230]), .op(N246_t0) );
fim FAN_N246_1 ( .fault(fault), .net(N246), .FEN(FEN[231]), .op(N246_t1) );
fim FAN_N246_2 ( .fault(fault), .net(N246), .FEN(FEN[232]), .op(N246_t2) );
fim FAN_N246_3 ( .fault(fault), .net(N246), .FEN(FEN[233]), .op(N246_t3) );
fim FAN_N246_4 ( .fault(fault), .net(N246), .FEN(FEN[234]), .op(N246_t4) );
fim FAN_N246_5 ( .fault(fault), .net(N246), .FEN(FEN[235]), .op(N246_t5) );
fim FAN_N11_0 ( .fault(fault), .net(N11), .FEN(FEN[236]), .op(N11_t0) );
fim FAN_N11_1 ( .fault(fault), .net(N11), .FEN(FEN[237]), .op(N11_t1) );
fim FAN_N256_0 ( .fault(fault), .net(N256), .FEN(FEN[238]), .op(N256_t0) );
fim FAN_N256_1 ( .fault(fault), .net(N256), .FEN(FEN[239]), .op(N256_t1) );
fim FAN_N259_0 ( .fault(fault), .net(N259), .FEN(FEN[240]), .op(N259_t0) );
fim FAN_N259_1 ( .fault(fault), .net(N259), .FEN(FEN[241]), .op(N259_t1) );
fim FAN_N319_0 ( .fault(fault), .net(N319), .FEN(FEN[242]), .op(N319_t0) );
fim FAN_N319_1 ( .fault(fault), .net(N319), .FEN(FEN[243]), .op(N319_t1) );
fim FAN_N322_0 ( .fault(fault), .net(N322), .FEN(FEN[244]), .op(N322_t0) );
fim FAN_N322_1 ( .fault(fault), .net(N322), .FEN(FEN[245]), .op(N322_t1) );
fim FAN_N328_0 ( .fault(fault), .net(N328), .FEN(FEN[246]), .op(N328_t0) );
fim FAN_N328_1 ( .fault(fault), .net(N328), .FEN(FEN[247]), .op(N328_t1) );
fim FAN_N331_0 ( .fault(fault), .net(N331), .FEN(FEN[248]), .op(N331_t0) );
fim FAN_N331_1 ( .fault(fault), .net(N331), .FEN(FEN[249]), .op(N331_t1) );
fim FAN_N334_0 ( .fault(fault), .net(N334), .FEN(FEN[250]), .op(N334_t0) );
fim FAN_N334_1 ( .fault(fault), .net(N334), .FEN(FEN[251]), .op(N334_t1) );
fim FAN_N337_0 ( .fault(fault), .net(N337), .FEN(FEN[252]), .op(N337_t0) );
fim FAN_N337_1 ( .fault(fault), .net(N337), .FEN(FEN[253]), .op(N337_t1) );
fim FAN_N340_0 ( .fault(fault), .net(N340), .FEN(FEN[254]), .op(N340_t0) );
fim FAN_N340_1 ( .fault(fault), .net(N340), .FEN(FEN[255]), .op(N340_t1) );
fim FAN_N343_0 ( .fault(fault), .net(N343), .FEN(FEN[256]), .op(N343_t0) );
fim FAN_N343_1 ( .fault(fault), .net(N343), .FEN(FEN[257]), .op(N343_t1) );
fim FAN_N352_0 ( .fault(fault), .net(N352), .FEN(FEN[258]), .op(N352_t0) );
fim FAN_N352_1 ( .fault(fault), .net(N352), .FEN(FEN[259]), .op(N352_t1) );
fim FAN_N16_0 ( .fault(fault), .net(N16), .FEN(FEN[260]), .op(N16_t0) );
fim FAN_N16_1 ( .fault(fault), .net(N16), .FEN(FEN[261]), .op(N16_t1) );
fim FAN_N355_0 ( .fault(fault), .net(N355), .FEN(FEN[262]), .op(N355_t0) );
fim FAN_N355_1 ( .fault(fault), .net(N355), .FEN(FEN[263]), .op(N355_t1) );
fim FAN_N263_0 ( .fault(fault), .net(N263), .FEN(FEN[264]), .op(N263_t0) );
fim FAN_N263_1 ( .fault(fault), .net(N263), .FEN(FEN[265]), .op(N263_t1) );
fim FAN_N266_0 ( .fault(fault), .net(N266), .FEN(FEN[266]), .op(N266_t0) );
fim FAN_N266_1 ( .fault(fault), .net(N266), .FEN(FEN[267]), .op(N266_t1) );
fim FAN_N269_0 ( .fault(fault), .net(N269), .FEN(FEN[268]), .op(N269_t0) );
fim FAN_N269_1 ( .fault(fault), .net(N269), .FEN(FEN[269]), .op(N269_t1) );
fim FAN_N272_0 ( .fault(fault), .net(N272), .FEN(FEN[270]), .op(N272_t0) );
fim FAN_N272_1 ( .fault(fault), .net(N272), .FEN(FEN[271]), .op(N272_t1) );
fim FAN_N275_0 ( .fault(fault), .net(N275), .FEN(FEN[272]), .op(N275_t0) );
fim FAN_N275_1 ( .fault(fault), .net(N275), .FEN(FEN[273]), .op(N275_t1) );
fim FAN_N278_0 ( .fault(fault), .net(N278), .FEN(FEN[274]), .op(N278_t0) );
fim FAN_N278_1 ( .fault(fault), .net(N278), .FEN(FEN[275]), .op(N278_t1) );
fim FAN_N281_0 ( .fault(fault), .net(N281), .FEN(FEN[276]), .op(N281_t0) );
fim FAN_N281_1 ( .fault(fault), .net(N281), .FEN(FEN[277]), .op(N281_t1) );
fim FAN_N284_0 ( .fault(fault), .net(N284), .FEN(FEN[278]), .op(N284_t0) );
fim FAN_N284_1 ( .fault(fault), .net(N284), .FEN(FEN[279]), .op(N284_t1) );
fim FAN_N287_0 ( .fault(fault), .net(N287), .FEN(FEN[280]), .op(N287_t0) );
fim FAN_N287_1 ( .fault(fault), .net(N287), .FEN(FEN[281]), .op(N287_t1) );
fim FAN_N29_0 ( .fault(fault), .net(N29), .FEN(FEN[282]), .op(N29_t0) );
fim FAN_N29_1 ( .fault(fault), .net(N29), .FEN(FEN[283]), .op(N29_t1) );
fim FAN_N294_0 ( .fault(fault), .net(N294), .FEN(FEN[284]), .op(N294_t0) );
fim FAN_N294_1 ( .fault(fault), .net(N294), .FEN(FEN[285]), .op(N294_t1) );
fim FAN_N313_0 ( .fault(fault), .net(N313), .FEN(FEN[286]), .op(N313_t0) );
fim FAN_N313_1 ( .fault(fault), .net(N313), .FEN(FEN[287]), .op(N313_t1) );
fim FAN_N316_0 ( .fault(fault), .net(N316), .FEN(FEN[288]), .op(N316_t0) );
fim FAN_N316_1 ( .fault(fault), .net(N316), .FEN(FEN[289]), .op(N316_t1) );
fim FAN_N346_0 ( .fault(fault), .net(N346), .FEN(FEN[290]), .op(N346_t0) );
fim FAN_N346_1 ( .fault(fault), .net(N346), .FEN(FEN[291]), .op(N346_t1) );
fim FAN_N349_0 ( .fault(fault), .net(N349), .FEN(FEN[292]), .op(N349_t0) );
fim FAN_N349_1 ( .fault(fault), .net(N349), .FEN(FEN[293]), .op(N349_t1) );
fim FAN_N500_0 ( .fault(fault), .net(N500), .FEN(FEN[294]), .op(N500_t0) );
fim FAN_N500_1 ( .fault(fault), .net(N500), .FEN(FEN[295]), .op(N500_t1) );
fim FAN_N325_0 ( .fault(fault), .net(N325), .FEN(FEN[296]), .op(N325_t0) );
fim FAN_N325_1 ( .fault(fault), .net(N325), .FEN(FEN[297]), .op(N325_t1) );
fim FAN_N651_0 ( .fault(fault), .net(N651), .FEN(FEN[298]), .op(N651_t0) );
fim FAN_N651_1 ( .fault(fault), .net(N651), .FEN(FEN[299]), .op(N651_t1) );
fim FAN_N651_2 ( .fault(fault), .net(N651), .FEN(FEN[300]), .op(N651_t2) );
fim FAN_N231_0 ( .fault(fault), .net(N231), .FEN(FEN[301]), .op(N231_t0) );
fim FAN_N231_1 ( .fault(fault), .net(N231), .FEN(FEN[302]), .op(N231_t1) );
fim FAN_N544_0 ( .fault(fault), .net(N544), .FEN(FEN[303]), .op(N544_t0) );
fim FAN_N544_1 ( .fault(fault), .net(N544), .FEN(FEN[304]), .op(N544_t1) );
fim FAN_N547_0 ( .fault(fault), .net(N547), .FEN(FEN[305]), .op(N547_t0) );
fim FAN_N547_1 ( .fault(fault), .net(N547), .FEN(FEN[306]), .op(N547_t1) );
fim FAN_N503_0 ( .fault(fault), .net(N503), .FEN(FEN[307]), .op(N503_t0) );
fim FAN_N503_1 ( .fault(fault), .net(N503), .FEN(FEN[308]), .op(N503_t1) );
fim FAN_N509_0 ( .fault(fault), .net(N509), .FEN(FEN[309]), .op(N509_t0) );
fim FAN_N509_1 ( .fault(fault), .net(N509), .FEN(FEN[310]), .op(N509_t1) );
fim FAN_N509_2 ( .fault(fault), .net(N509), .FEN(FEN[311]), .op(N509_t2) );
fim FAN_N509_3 ( .fault(fault), .net(N509), .FEN(FEN[312]), .op(N509_t3) );
fim FAN_N509_4 ( .fault(fault), .net(N509), .FEN(FEN[313]), .op(N509_t4) );
fim FAN_N509_5 ( .fault(fault), .net(N509), .FEN(FEN[314]), .op(N509_t5) );
fim FAN_N509_6 ( .fault(fault), .net(N509), .FEN(FEN[315]), .op(N509_t6) );
fim FAN_N509_7 ( .fault(fault), .net(N509), .FEN(FEN[316]), .op(N509_t7) );
fim FAN_N509_8 ( .fault(fault), .net(N509), .FEN(FEN[317]), .op(N509_t8) );
fim FAN_N509_9 ( .fault(fault), .net(N509), .FEN(FEN[318]), .op(N509_t9) );
fim FAN_N509_10 ( .fault(fault), .net(N509), .FEN(FEN[319]), .op(N509_t10) );
fim FAN_N521_0 ( .fault(fault), .net(N521), .FEN(FEN[320]), .op(N521_t0) );
fim FAN_N521_1 ( .fault(fault), .net(N521), .FEN(FEN[321]), .op(N521_t1) );
fim FAN_N521_2 ( .fault(fault), .net(N521), .FEN(FEN[322]), .op(N521_t2) );
fim FAN_N521_3 ( .fault(fault), .net(N521), .FEN(FEN[323]), .op(N521_t3) );
fim FAN_N521_4 ( .fault(fault), .net(N521), .FEN(FEN[324]), .op(N521_t4) );
fim FAN_N521_5 ( .fault(fault), .net(N521), .FEN(FEN[325]), .op(N521_t5) );
fim FAN_N521_6 ( .fault(fault), .net(N521), .FEN(FEN[326]), .op(N521_t6) );
fim FAN_N521_7 ( .fault(fault), .net(N521), .FEN(FEN[327]), .op(N521_t7) );
fim FAN_N521_8 ( .fault(fault), .net(N521), .FEN(FEN[328]), .op(N521_t8) );
fim FAN_N521_9 ( .fault(fault), .net(N521), .FEN(FEN[329]), .op(N521_t9) );
fim FAN_N521_10 ( .fault(fault), .net(N521), .FEN(FEN[330]), .op(N521_t10) );
fim FAN_N537_0 ( .fault(fault), .net(N537), .FEN(FEN[331]), .op(N537_t0) );
fim FAN_N537_1 ( .fault(fault), .net(N537), .FEN(FEN[332]), .op(N537_t1) );
fim FAN_N537_2 ( .fault(fault), .net(N537), .FEN(FEN[333]), .op(N537_t2) );
fim FAN_N537_3 ( .fault(fault), .net(N537), .FEN(FEN[334]), .op(N537_t3) );
fim FAN_N537_4 ( .fault(fault), .net(N537), .FEN(FEN[335]), .op(N537_t4) );
fim FAN_N550_0 ( .fault(fault), .net(N550), .FEN(FEN[336]), .op(N550_t0) );
fim FAN_N550_1 ( .fault(fault), .net(N550), .FEN(FEN[337]), .op(N550_t1) );
fim FAN_N550_2 ( .fault(fault), .net(N550), .FEN(FEN[338]), .op(N550_t2) );
fim FAN_N550_3 ( .fault(fault), .net(N550), .FEN(FEN[339]), .op(N550_t3) );
fim FAN_N550_4 ( .fault(fault), .net(N550), .FEN(FEN[340]), .op(N550_t4) );
fim FAN_N550_5 ( .fault(fault), .net(N550), .FEN(FEN[341]), .op(N550_t5) );
fim FAN_N550_6 ( .fault(fault), .net(N550), .FEN(FEN[342]), .op(N550_t6) );
fim FAN_N550_7 ( .fault(fault), .net(N550), .FEN(FEN[343]), .op(N550_t7) );
fim FAN_N550_8 ( .fault(fault), .net(N550), .FEN(FEN[344]), .op(N550_t8) );
fim FAN_N550_9 ( .fault(fault), .net(N550), .FEN(FEN[345]), .op(N550_t9) );
fim FAN_N550_10 ( .fault(fault), .net(N550), .FEN(FEN[346]), .op(N550_t10) );
fim FAN_N562_0 ( .fault(fault), .net(N562), .FEN(FEN[347]), .op(N562_t0) );
fim FAN_N562_1 ( .fault(fault), .net(N562), .FEN(FEN[348]), .op(N562_t1) );
fim FAN_N562_2 ( .fault(fault), .net(N562), .FEN(FEN[349]), .op(N562_t2) );
fim FAN_N562_3 ( .fault(fault), .net(N562), .FEN(FEN[350]), .op(N562_t3) );
fim FAN_N562_4 ( .fault(fault), .net(N562), .FEN(FEN[351]), .op(N562_t4) );
fim FAN_N562_5 ( .fault(fault), .net(N562), .FEN(FEN[352]), .op(N562_t5) );
fim FAN_N562_6 ( .fault(fault), .net(N562), .FEN(FEN[353]), .op(N562_t6) );
fim FAN_N562_7 ( .fault(fault), .net(N562), .FEN(FEN[354]), .op(N562_t7) );
fim FAN_N562_8 ( .fault(fault), .net(N562), .FEN(FEN[355]), .op(N562_t8) );
fim FAN_N562_9 ( .fault(fault), .net(N562), .FEN(FEN[356]), .op(N562_t9) );
fim FAN_N562_10 ( .fault(fault), .net(N562), .FEN(FEN[357]), .op(N562_t10) );
fim FAN_N582_0 ( .fault(fault), .net(N582), .FEN(FEN[358]), .op(N582_t0) );
fim FAN_N582_1 ( .fault(fault), .net(N582), .FEN(FEN[359]), .op(N582_t1) );
fim FAN_N582_2 ( .fault(fault), .net(N582), .FEN(FEN[360]), .op(N582_t2) );
fim FAN_N582_3 ( .fault(fault), .net(N582), .FEN(FEN[361]), .op(N582_t3) );
fim FAN_N582_4 ( .fault(fault), .net(N582), .FEN(FEN[362]), .op(N582_t4) );
fim FAN_N582_5 ( .fault(fault), .net(N582), .FEN(FEN[363]), .op(N582_t5) );
fim FAN_N582_6 ( .fault(fault), .net(N582), .FEN(FEN[364]), .op(N582_t6) );
fim FAN_N582_7 ( .fault(fault), .net(N582), .FEN(FEN[365]), .op(N582_t7) );
fim FAN_N582_8 ( .fault(fault), .net(N582), .FEN(FEN[366]), .op(N582_t8) );
fim FAN_N582_9 ( .fault(fault), .net(N582), .FEN(FEN[367]), .op(N582_t9) );
fim FAN_N582_10 ( .fault(fault), .net(N582), .FEN(FEN[368]), .op(N582_t10) );
fim FAN_N594_0 ( .fault(fault), .net(N594), .FEN(FEN[369]), .op(N594_t0) );
fim FAN_N594_1 ( .fault(fault), .net(N594), .FEN(FEN[370]), .op(N594_t1) );
fim FAN_N594_2 ( .fault(fault), .net(N594), .FEN(FEN[371]), .op(N594_t2) );
fim FAN_N594_3 ( .fault(fault), .net(N594), .FEN(FEN[372]), .op(N594_t3) );
fim FAN_N594_4 ( .fault(fault), .net(N594), .FEN(FEN[373]), .op(N594_t4) );
fim FAN_N594_5 ( .fault(fault), .net(N594), .FEN(FEN[374]), .op(N594_t5) );
fim FAN_N594_6 ( .fault(fault), .net(N594), .FEN(FEN[375]), .op(N594_t6) );
fim FAN_N594_7 ( .fault(fault), .net(N594), .FEN(FEN[376]), .op(N594_t7) );
fim FAN_N594_8 ( .fault(fault), .net(N594), .FEN(FEN[377]), .op(N594_t8) );
fim FAN_N594_9 ( .fault(fault), .net(N594), .FEN(FEN[378]), .op(N594_t9) );
fim FAN_N594_10 ( .fault(fault), .net(N594), .FEN(FEN[379]), .op(N594_t10) );
fim FAN_N741_0 ( .fault(fault), .net(N741), .FEN(FEN[380]), .op(N741_t0) );
fim FAN_N741_1 ( .fault(fault), .net(N741), .FEN(FEN[381]), .op(N741_t1) );
fim FAN_N744_0 ( .fault(fault), .net(N744), .FEN(FEN[382]), .op(N744_t0) );
fim FAN_N744_1 ( .fault(fault), .net(N744), .FEN(FEN[383]), .op(N744_t1) );
fim FAN_N747_0 ( .fault(fault), .net(N747), .FEN(FEN[384]), .op(N747_t0) );
fim FAN_N747_1 ( .fault(fault), .net(N747), .FEN(FEN[385]), .op(N747_t1) );
fim FAN_N750_0 ( .fault(fault), .net(N750), .FEN(FEN[386]), .op(N750_t0) );
fim FAN_N750_1 ( .fault(fault), .net(N750), .FEN(FEN[387]), .op(N750_t1) );
fim FAN_N753_0 ( .fault(fault), .net(N753), .FEN(FEN[388]), .op(N753_t0) );
fim FAN_N753_1 ( .fault(fault), .net(N753), .FEN(FEN[389]), .op(N753_t1) );
fim FAN_N613_0 ( .fault(fault), .net(N613), .FEN(FEN[390]), .op(N613_t0) );
fim FAN_N613_1 ( .fault(fault), .net(N613), .FEN(FEN[391]), .op(N613_t1) );
fim FAN_N613_2 ( .fault(fault), .net(N613), .FEN(FEN[392]), .op(N613_t2) );
fim FAN_N613_3 ( .fault(fault), .net(N613), .FEN(FEN[393]), .op(N613_t3) );
fim FAN_N613_4 ( .fault(fault), .net(N613), .FEN(FEN[394]), .op(N613_t4) );
fim FAN_N613_5 ( .fault(fault), .net(N613), .FEN(FEN[395]), .op(N613_t5) );
fim FAN_N613_6 ( .fault(fault), .net(N613), .FEN(FEN[396]), .op(N613_t6) );
fim FAN_N613_7 ( .fault(fault), .net(N613), .FEN(FEN[397]), .op(N613_t7) );
fim FAN_N613_8 ( .fault(fault), .net(N613), .FEN(FEN[398]), .op(N613_t8) );
fim FAN_N613_9 ( .fault(fault), .net(N613), .FEN(FEN[399]), .op(N613_t9) );
fim FAN_N613_10 ( .fault(fault), .net(N613), .FEN(FEN[400]), .op(N613_t10) );
fim FAN_N625_0 ( .fault(fault), .net(N625), .FEN(FEN[401]), .op(N625_t0) );
fim FAN_N625_1 ( .fault(fault), .net(N625), .FEN(FEN[402]), .op(N625_t1) );
fim FAN_N625_2 ( .fault(fault), .net(N625), .FEN(FEN[403]), .op(N625_t2) );
fim FAN_N625_3 ( .fault(fault), .net(N625), .FEN(FEN[404]), .op(N625_t3) );
fim FAN_N625_4 ( .fault(fault), .net(N625), .FEN(FEN[405]), .op(N625_t4) );
fim FAN_N625_5 ( .fault(fault), .net(N625), .FEN(FEN[406]), .op(N625_t5) );
fim FAN_N625_6 ( .fault(fault), .net(N625), .FEN(FEN[407]), .op(N625_t6) );
fim FAN_N625_7 ( .fault(fault), .net(N625), .FEN(FEN[408]), .op(N625_t7) );
fim FAN_N625_8 ( .fault(fault), .net(N625), .FEN(FEN[409]), .op(N625_t8) );
fim FAN_N625_9 ( .fault(fault), .net(N625), .FEN(FEN[410]), .op(N625_t9) );
fim FAN_N625_10 ( .fault(fault), .net(N625), .FEN(FEN[411]), .op(N625_t10) );
fim FAN_N637_0 ( .fault(fault), .net(N637), .FEN(FEN[412]), .op(N637_t0) );
fim FAN_N637_1 ( .fault(fault), .net(N637), .FEN(FEN[413]), .op(N637_t1) );
fim FAN_N637_2 ( .fault(fault), .net(N637), .FEN(FEN[414]), .op(N637_t2) );
fim FAN_N637_3 ( .fault(fault), .net(N637), .FEN(FEN[415]), .op(N637_t3) );
fim FAN_N637_4 ( .fault(fault), .net(N637), .FEN(FEN[416]), .op(N637_t4) );
fim FAN_N643_0 ( .fault(fault), .net(N643), .FEN(FEN[417]), .op(N643_t0) );
fim FAN_N643_1 ( .fault(fault), .net(N643), .FEN(FEN[418]), .op(N643_t1) );
fim FAN_N643_2 ( .fault(fault), .net(N643), .FEN(FEN[419]), .op(N643_t2) );
fim FAN_N643_3 ( .fault(fault), .net(N643), .FEN(FEN[420]), .op(N643_t3) );
fim FAN_N643_4 ( .fault(fault), .net(N643), .FEN(FEN[421]), .op(N643_t4) );
fim FAN_N643_5 ( .fault(fault), .net(N643), .FEN(FEN[422]), .op(N643_t5) );
fim FAN_N768_0 ( .fault(fault), .net(N768), .FEN(FEN[423]), .op(N768_t0) );
fim FAN_N768_1 ( .fault(fault), .net(N768), .FEN(FEN[424]), .op(N768_t1) );
fim FAN_N771_0 ( .fault(fault), .net(N771), .FEN(FEN[425]), .op(N771_t0) );
fim FAN_N771_1 ( .fault(fault), .net(N771), .FEN(FEN[426]), .op(N771_t1) );
fim FAN_N774_0 ( .fault(fault), .net(N774), .FEN(FEN[427]), .op(N774_t0) );
fim FAN_N774_1 ( .fault(fault), .net(N774), .FEN(FEN[428]), .op(N774_t1) );
fim FAN_N777_0 ( .fault(fault), .net(N777), .FEN(FEN[429]), .op(N777_t0) );
fim FAN_N777_1 ( .fault(fault), .net(N777), .FEN(FEN[430]), .op(N777_t1) );
fim FAN_N780_0 ( .fault(fault), .net(N780), .FEN(FEN[431]), .op(N780_t0) );
fim FAN_N780_1 ( .fault(fault), .net(N780), .FEN(FEN[432]), .op(N780_t1) );
fim FAN_N506_0 ( .fault(fault), .net(N506), .FEN(FEN[433]), .op(N506_t0) );
fim FAN_N506_1 ( .fault(fault), .net(N506), .FEN(FEN[434]), .op(N506_t1) );
fim FAN_N693_0 ( .fault(fault), .net(N693), .FEN(FEN[435]), .op(N693_t0) );
fim FAN_N693_1 ( .fault(fault), .net(N693), .FEN(FEN[436]), .op(N693_t1) );
fim FAN_N693_2 ( .fault(fault), .net(N693), .FEN(FEN[437]), .op(N693_t2) );
fim FAN_N693_3 ( .fault(fault), .net(N693), .FEN(FEN[438]), .op(N693_t3) );
fim FAN_N693_4 ( .fault(fault), .net(N693), .FEN(FEN[439]), .op(N693_t4) );
fim FAN_N699_0 ( .fault(fault), .net(N699), .FEN(FEN[440]), .op(N699_t0) );
fim FAN_N699_1 ( .fault(fault), .net(N699), .FEN(FEN[441]), .op(N699_t1) );
fim FAN_N699_2 ( .fault(fault), .net(N699), .FEN(FEN[442]), .op(N699_t2) );
fim FAN_N699_3 ( .fault(fault), .net(N699), .FEN(FEN[443]), .op(N699_t3) );
fim FAN_N699_4 ( .fault(fault), .net(N699), .FEN(FEN[444]), .op(N699_t4) );
fim FAN_N735_0 ( .fault(fault), .net(N735), .FEN(FEN[445]), .op(N735_t0) );
fim FAN_N735_1 ( .fault(fault), .net(N735), .FEN(FEN[446]), .op(N735_t1) );
fim FAN_N738_0 ( .fault(fault), .net(N738), .FEN(FEN[447]), .op(N738_t0) );
fim FAN_N738_1 ( .fault(fault), .net(N738), .FEN(FEN[448]), .op(N738_t1) );
fim FAN_N756_0 ( .fault(fault), .net(N756), .FEN(FEN[449]), .op(N756_t0) );
fim FAN_N756_1 ( .fault(fault), .net(N756), .FEN(FEN[450]), .op(N756_t1) );
fim FAN_N759_0 ( .fault(fault), .net(N759), .FEN(FEN[451]), .op(N759_t0) );
fim FAN_N759_1 ( .fault(fault), .net(N759), .FEN(FEN[452]), .op(N759_t1) );
fim FAN_N762_0 ( .fault(fault), .net(N762), .FEN(FEN[453]), .op(N762_t0) );
fim FAN_N762_1 ( .fault(fault), .net(N762), .FEN(FEN[454]), .op(N762_t1) );
fim FAN_N765_0 ( .fault(fault), .net(N765), .FEN(FEN[455]), .op(N765_t0) );
fim FAN_N765_1 ( .fault(fault), .net(N765), .FEN(FEN[456]), .op(N765_t1) );
fim FAN_N574_0 ( .fault(fault), .net(N574), .FEN(FEN[457]), .op(N574_t0) );
fim FAN_N574_1 ( .fault(fault), .net(N574), .FEN(FEN[458]), .op(N574_t1) );
fim FAN_N574_2 ( .fault(fault), .net(N574), .FEN(FEN[459]), .op(N574_t2) );
fim FAN_N578_0 ( .fault(fault), .net(N578), .FEN(FEN[460]), .op(N578_t0) );
fim FAN_N578_1 ( .fault(fault), .net(N578), .FEN(FEN[461]), .op(N578_t1) );
fim FAN_N578_2 ( .fault(fault), .net(N578), .FEN(FEN[462]), .op(N578_t2) );
fim FAN_N655_0 ( .fault(fault), .net(N655), .FEN(FEN[463]), .op(N655_t0) );
fim FAN_N655_1 ( .fault(fault), .net(N655), .FEN(FEN[464]), .op(N655_t1) );
fim FAN_N655_2 ( .fault(fault), .net(N655), .FEN(FEN[465]), .op(N655_t2) );
fim FAN_N659_0 ( .fault(fault), .net(N659), .FEN(FEN[466]), .op(N659_t0) );
fim FAN_N659_1 ( .fault(fault), .net(N659), .FEN(FEN[467]), .op(N659_t1) );
fim FAN_N659_2 ( .fault(fault), .net(N659), .FEN(FEN[468]), .op(N659_t2) );
fim FAN_N663_0 ( .fault(fault), .net(N663), .FEN(FEN[469]), .op(N663_t0) );
fim FAN_N663_1 ( .fault(fault), .net(N663), .FEN(FEN[470]), .op(N663_t1) );
fim FAN_N663_2 ( .fault(fault), .net(N663), .FEN(FEN[471]), .op(N663_t2) );
fim FAN_N667_0 ( .fault(fault), .net(N667), .FEN(FEN[472]), .op(N667_t0) );
fim FAN_N667_1 ( .fault(fault), .net(N667), .FEN(FEN[473]), .op(N667_t1) );
fim FAN_N667_2 ( .fault(fault), .net(N667), .FEN(FEN[474]), .op(N667_t2) );
fim FAN_N671_0 ( .fault(fault), .net(N671), .FEN(FEN[475]), .op(N671_t0) );
fim FAN_N671_1 ( .fault(fault), .net(N671), .FEN(FEN[476]), .op(N671_t1) );
fim FAN_N671_2 ( .fault(fault), .net(N671), .FEN(FEN[477]), .op(N671_t2) );
fim FAN_N675_0 ( .fault(fault), .net(N675), .FEN(FEN[478]), .op(N675_t0) );
fim FAN_N675_1 ( .fault(fault), .net(N675), .FEN(FEN[479]), .op(N675_t1) );
fim FAN_N675_2 ( .fault(fault), .net(N675), .FEN(FEN[480]), .op(N675_t2) );
fim FAN_N679_0 ( .fault(fault), .net(N679), .FEN(FEN[481]), .op(N679_t0) );
fim FAN_N679_1 ( .fault(fault), .net(N679), .FEN(FEN[482]), .op(N679_t1) );
fim FAN_N679_2 ( .fault(fault), .net(N679), .FEN(FEN[483]), .op(N679_t2) );
fim FAN_N683_0 ( .fault(fault), .net(N683), .FEN(FEN[484]), .op(N683_t0) );
fim FAN_N683_1 ( .fault(fault), .net(N683), .FEN(FEN[485]), .op(N683_t1) );
fim FAN_N683_2 ( .fault(fault), .net(N683), .FEN(FEN[486]), .op(N683_t2) );
fim FAN_N783_0 ( .fault(fault), .net(N783), .FEN(FEN[487]), .op(N783_t0) );
fim FAN_N783_1 ( .fault(fault), .net(N783), .FEN(FEN[488]), .op(N783_t1) );
fim FAN_N786_0 ( .fault(fault), .net(N786), .FEN(FEN[489]), .op(N786_t0) );
fim FAN_N786_1 ( .fault(fault), .net(N786), .FEN(FEN[490]), .op(N786_t1) );
fim FAN_N687_0 ( .fault(fault), .net(N687), .FEN(FEN[491]), .op(N687_t0) );
fim FAN_N687_1 ( .fault(fault), .net(N687), .FEN(FEN[492]), .op(N687_t1) );
fim FAN_N687_2 ( .fault(fault), .net(N687), .FEN(FEN[493]), .op(N687_t2) );
fim FAN_N687_3 ( .fault(fault), .net(N687), .FEN(FEN[494]), .op(N687_t3) );
fim FAN_N687_4 ( .fault(fault), .net(N687), .FEN(FEN[495]), .op(N687_t4) );
fim FAN_N705_0 ( .fault(fault), .net(N705), .FEN(FEN[496]), .op(N705_t0) );
fim FAN_N705_1 ( .fault(fault), .net(N705), .FEN(FEN[497]), .op(N705_t1) );
fim FAN_N705_2 ( .fault(fault), .net(N705), .FEN(FEN[498]), .op(N705_t2) );
fim FAN_N705_3 ( .fault(fault), .net(N705), .FEN(FEN[499]), .op(N705_t3) );
fim FAN_N705_4 ( .fault(fault), .net(N705), .FEN(FEN[500]), .op(N705_t4) );
fim FAN_N711_0 ( .fault(fault), .net(N711), .FEN(FEN[501]), .op(N711_t0) );
fim FAN_N711_1 ( .fault(fault), .net(N711), .FEN(FEN[502]), .op(N711_t1) );
fim FAN_N711_2 ( .fault(fault), .net(N711), .FEN(FEN[503]), .op(N711_t2) );
fim FAN_N715_0 ( .fault(fault), .net(N715), .FEN(FEN[504]), .op(N715_t0) );
fim FAN_N715_1 ( .fault(fault), .net(N715), .FEN(FEN[505]), .op(N715_t1) );
fim FAN_N715_2 ( .fault(fault), .net(N715), .FEN(FEN[506]), .op(N715_t2) );
fim FAN_N719_0 ( .fault(fault), .net(N719), .FEN(FEN[507]), .op(N719_t0) );
fim FAN_N719_1 ( .fault(fault), .net(N719), .FEN(FEN[508]), .op(N719_t1) );
fim FAN_N719_2 ( .fault(fault), .net(N719), .FEN(FEN[509]), .op(N719_t2) );
fim FAN_N723_0 ( .fault(fault), .net(N723), .FEN(FEN[510]), .op(N723_t0) );
fim FAN_N723_1 ( .fault(fault), .net(N723), .FEN(FEN[511]), .op(N723_t1) );
fim FAN_N723_2 ( .fault(fault), .net(N723), .FEN(FEN[512]), .op(N723_t2) );
fim FAN_N1034_0 ( .fault(fault), .net(N1034), .FEN(FEN[513]), .op(N1034_t0) );
fim FAN_N1034_1 ( .fault(fault), .net(N1034), .FEN(FEN[514]), .op(N1034_t1) );
fim FAN_N1042_0 ( .fault(fault), .net(N1042), .FEN(FEN[515]), .op(N1042_t0) );
fim FAN_N1042_1 ( .fault(fault), .net(N1042), .FEN(FEN[516]), .op(N1042_t1) );
fim FAN_N1042_2 ( .fault(fault), .net(N1042), .FEN(FEN[517]), .op(N1042_t2) );
fim FAN_N1042_3 ( .fault(fault), .net(N1042), .FEN(FEN[518]), .op(N1042_t3) );
fim FAN_N1042_4 ( .fault(fault), .net(N1042), .FEN(FEN[519]), .op(N1042_t4) );
fim FAN_N1042_5 ( .fault(fault), .net(N1042), .FEN(FEN[520]), .op(N1042_t5) );
fim FAN_N1042_6 ( .fault(fault), .net(N1042), .FEN(FEN[521]), .op(N1042_t6) );
fim FAN_N1042_7 ( .fault(fault), .net(N1042), .FEN(FEN[522]), .op(N1042_t7) );
fim FAN_N1042_8 ( .fault(fault), .net(N1042), .FEN(FEN[523]), .op(N1042_t8) );
fim FAN_N1042_9 ( .fault(fault), .net(N1042), .FEN(FEN[524]), .op(N1042_t9) );
fim FAN_N1053_0 ( .fault(fault), .net(N1053), .FEN(FEN[525]), .op(N1053_t0) );
fim FAN_N1053_1 ( .fault(fault), .net(N1053), .FEN(FEN[526]), .op(N1053_t1) );
fim FAN_N1053_2 ( .fault(fault), .net(N1053), .FEN(FEN[527]), .op(N1053_t2) );
fim FAN_N1053_3 ( .fault(fault), .net(N1053), .FEN(FEN[528]), .op(N1053_t3) );
fim FAN_N1053_4 ( .fault(fault), .net(N1053), .FEN(FEN[529]), .op(N1053_t4) );
fim FAN_N1053_5 ( .fault(fault), .net(N1053), .FEN(FEN[530]), .op(N1053_t5) );
fim FAN_N1053_6 ( .fault(fault), .net(N1053), .FEN(FEN[531]), .op(N1053_t6) );
fim FAN_N1053_7 ( .fault(fault), .net(N1053), .FEN(FEN[532]), .op(N1053_t7) );
fim FAN_N1053_8 ( .fault(fault), .net(N1053), .FEN(FEN[533]), .op(N1053_t8) );
fim FAN_N1053_9 ( .fault(fault), .net(N1053), .FEN(FEN[534]), .op(N1053_t9) );
fim FAN_N1075_0 ( .fault(fault), .net(N1075), .FEN(FEN[535]), .op(N1075_t0) );
fim FAN_N1075_1 ( .fault(fault), .net(N1075), .FEN(FEN[536]), .op(N1075_t1) );
fim FAN_N1075_2 ( .fault(fault), .net(N1075), .FEN(FEN[537]), .op(N1075_t2) );
fim FAN_N1075_3 ( .fault(fault), .net(N1075), .FEN(FEN[538]), .op(N1075_t3) );
fim FAN_N1075_4 ( .fault(fault), .net(N1075), .FEN(FEN[539]), .op(N1075_t4) );
fim FAN_N1075_5 ( .fault(fault), .net(N1075), .FEN(FEN[540]), .op(N1075_t5) );
fim FAN_N1075_6 ( .fault(fault), .net(N1075), .FEN(FEN[541]), .op(N1075_t6) );
fim FAN_N1075_7 ( .fault(fault), .net(N1075), .FEN(FEN[542]), .op(N1075_t7) );
fim FAN_N1075_8 ( .fault(fault), .net(N1075), .FEN(FEN[543]), .op(N1075_t8) );
fim FAN_N1075_9 ( .fault(fault), .net(N1075), .FEN(FEN[544]), .op(N1075_t9) );
fim FAN_N1086_0 ( .fault(fault), .net(N1086), .FEN(FEN[545]), .op(N1086_t0) );
fim FAN_N1086_1 ( .fault(fault), .net(N1086), .FEN(FEN[546]), .op(N1086_t1) );
fim FAN_N1086_2 ( .fault(fault), .net(N1086), .FEN(FEN[547]), .op(N1086_t2) );
fim FAN_N1086_3 ( .fault(fault), .net(N1086), .FEN(FEN[548]), .op(N1086_t3) );
fim FAN_N1086_4 ( .fault(fault), .net(N1086), .FEN(FEN[549]), .op(N1086_t4) );
fim FAN_N1086_5 ( .fault(fault), .net(N1086), .FEN(FEN[550]), .op(N1086_t5) );
fim FAN_N1086_6 ( .fault(fault), .net(N1086), .FEN(FEN[551]), .op(N1086_t6) );
fim FAN_N1086_7 ( .fault(fault), .net(N1086), .FEN(FEN[552]), .op(N1086_t7) );
fim FAN_N1086_8 ( .fault(fault), .net(N1086), .FEN(FEN[553]), .op(N1086_t8) );
fim FAN_N1086_9 ( .fault(fault), .net(N1086), .FEN(FEN[554]), .op(N1086_t9) );
fim FAN_N1102_0 ( .fault(fault), .net(N1102), .FEN(FEN[555]), .op(N1102_t0) );
fim FAN_N1102_1 ( .fault(fault), .net(N1102), .FEN(FEN[556]), .op(N1102_t1) );
fim FAN_N1102_2 ( .fault(fault), .net(N1102), .FEN(FEN[557]), .op(N1102_t2) );
fim FAN_N1102_3 ( .fault(fault), .net(N1102), .FEN(FEN[558]), .op(N1102_t3) );
fim FAN_N1102_4 ( .fault(fault), .net(N1102), .FEN(FEN[559]), .op(N1102_t4) );
fim FAN_N1102_5 ( .fault(fault), .net(N1102), .FEN(FEN[560]), .op(N1102_t5) );
fim FAN_N1102_6 ( .fault(fault), .net(N1102), .FEN(FEN[561]), .op(N1102_t6) );
fim FAN_N1102_7 ( .fault(fault), .net(N1102), .FEN(FEN[562]), .op(N1102_t7) );
fim FAN_N1102_8 ( .fault(fault), .net(N1102), .FEN(FEN[563]), .op(N1102_t8) );
fim FAN_N1102_9 ( .fault(fault), .net(N1102), .FEN(FEN[564]), .op(N1102_t9) );
fim FAN_N1113_0 ( .fault(fault), .net(N1113), .FEN(FEN[565]), .op(N1113_t0) );
fim FAN_N1113_1 ( .fault(fault), .net(N1113), .FEN(FEN[566]), .op(N1113_t1) );
fim FAN_N1113_2 ( .fault(fault), .net(N1113), .FEN(FEN[567]), .op(N1113_t2) );
fim FAN_N1113_3 ( .fault(fault), .net(N1113), .FEN(FEN[568]), .op(N1113_t3) );
fim FAN_N1113_4 ( .fault(fault), .net(N1113), .FEN(FEN[569]), .op(N1113_t4) );
fim FAN_N1113_5 ( .fault(fault), .net(N1113), .FEN(FEN[570]), .op(N1113_t5) );
fim FAN_N1113_6 ( .fault(fault), .net(N1113), .FEN(FEN[571]), .op(N1113_t6) );
fim FAN_N1113_7 ( .fault(fault), .net(N1113), .FEN(FEN[572]), .op(N1113_t7) );
fim FAN_N1113_8 ( .fault(fault), .net(N1113), .FEN(FEN[573]), .op(N1113_t8) );
fim FAN_N1113_9 ( .fault(fault), .net(N1113), .FEN(FEN[574]), .op(N1113_t9) );
fim FAN_N1129_0 ( .fault(fault), .net(N1129), .FEN(FEN[575]), .op(N1129_t0) );
fim FAN_N1129_1 ( .fault(fault), .net(N1129), .FEN(FEN[576]), .op(N1129_t1) );
fim FAN_N1129_2 ( .fault(fault), .net(N1129), .FEN(FEN[577]), .op(N1129_t2) );
fim FAN_N1133_0 ( .fault(fault), .net(N1133), .FEN(FEN[578]), .op(N1133_t0) );
fim FAN_N1133_1 ( .fault(fault), .net(N1133), .FEN(FEN[579]), .op(N1133_t1) );
fim FAN_N1133_2 ( .fault(fault), .net(N1133), .FEN(FEN[580]), .op(N1133_t2) );
fim FAN_N1137_0 ( .fault(fault), .net(N1137), .FEN(FEN[581]), .op(N1137_t0) );
fim FAN_N1137_1 ( .fault(fault), .net(N1137), .FEN(FEN[582]), .op(N1137_t1) );
fim FAN_N1219_0 ( .fault(fault), .net(N1219), .FEN(FEN[583]), .op(N1219_t0) );
fim FAN_N1219_1 ( .fault(fault), .net(N1219), .FEN(FEN[584]), .op(N1219_t1) );
fim FAN_N1222_0 ( .fault(fault), .net(N1222), .FEN(FEN[585]), .op(N1222_t0) );
fim FAN_N1222_1 ( .fault(fault), .net(N1222), .FEN(FEN[586]), .op(N1222_t1) );
fim FAN_N1225_0 ( .fault(fault), .net(N1225), .FEN(FEN[587]), .op(N1225_t0) );
fim FAN_N1225_1 ( .fault(fault), .net(N1225), .FEN(FEN[588]), .op(N1225_t1) );
fim FAN_N1228_0 ( .fault(fault), .net(N1228), .FEN(FEN[589]), .op(N1228_t0) );
fim FAN_N1228_1 ( .fault(fault), .net(N1228), .FEN(FEN[590]), .op(N1228_t1) );
fim FAN_N1231_0 ( .fault(fault), .net(N1231), .FEN(FEN[591]), .op(N1231_t0) );
fim FAN_N1231_1 ( .fault(fault), .net(N1231), .FEN(FEN[592]), .op(N1231_t1) );
fim FAN_N1234_0 ( .fault(fault), .net(N1234), .FEN(FEN[593]), .op(N1234_t0) );
fim FAN_N1234_1 ( .fault(fault), .net(N1234), .FEN(FEN[594]), .op(N1234_t1) );
fim FAN_N1237_0 ( .fault(fault), .net(N1237), .FEN(FEN[595]), .op(N1237_t0) );
fim FAN_N1237_1 ( .fault(fault), .net(N1237), .FEN(FEN[596]), .op(N1237_t1) );
fim FAN_N1240_0 ( .fault(fault), .net(N1240), .FEN(FEN[597]), .op(N1240_t0) );
fim FAN_N1240_1 ( .fault(fault), .net(N1240), .FEN(FEN[598]), .op(N1240_t1) );
fim FAN_N1243_0 ( .fault(fault), .net(N1243), .FEN(FEN[599]), .op(N1243_t0) );
fim FAN_N1243_1 ( .fault(fault), .net(N1243), .FEN(FEN[600]), .op(N1243_t1) );
fim FAN_N1246_0 ( .fault(fault), .net(N1246), .FEN(FEN[601]), .op(N1246_t0) );
fim FAN_N1246_1 ( .fault(fault), .net(N1246), .FEN(FEN[602]), .op(N1246_t1) );
fim FAN_N1146_0 ( .fault(fault), .net(N1146), .FEN(FEN[603]), .op(N1146_t0) );
fim FAN_N1146_1 ( .fault(fault), .net(N1146), .FEN(FEN[604]), .op(N1146_t1) );
fim FAN_N1146_2 ( .fault(fault), .net(N1146), .FEN(FEN[605]), .op(N1146_t2) );
fim FAN_N1146_3 ( .fault(fault), .net(N1146), .FEN(FEN[606]), .op(N1146_t3) );
fim FAN_N1146_4 ( .fault(fault), .net(N1146), .FEN(FEN[607]), .op(N1146_t4) );
fim FAN_N1146_5 ( .fault(fault), .net(N1146), .FEN(FEN[608]), .op(N1146_t5) );
fim FAN_N1146_6 ( .fault(fault), .net(N1146), .FEN(FEN[609]), .op(N1146_t6) );
fim FAN_N1146_7 ( .fault(fault), .net(N1146), .FEN(FEN[610]), .op(N1146_t7) );
fim FAN_N1146_8 ( .fault(fault), .net(N1146), .FEN(FEN[611]), .op(N1146_t8) );
fim FAN_N1146_9 ( .fault(fault), .net(N1146), .FEN(FEN[612]), .op(N1146_t9) );
fim FAN_N1157_0 ( .fault(fault), .net(N1157), .FEN(FEN[613]), .op(N1157_t0) );
fim FAN_N1157_1 ( .fault(fault), .net(N1157), .FEN(FEN[614]), .op(N1157_t1) );
fim FAN_N1157_2 ( .fault(fault), .net(N1157), .FEN(FEN[615]), .op(N1157_t2) );
fim FAN_N1157_3 ( .fault(fault), .net(N1157), .FEN(FEN[616]), .op(N1157_t3) );
fim FAN_N1157_4 ( .fault(fault), .net(N1157), .FEN(FEN[617]), .op(N1157_t4) );
fim FAN_N1157_5 ( .fault(fault), .net(N1157), .FEN(FEN[618]), .op(N1157_t5) );
fim FAN_N1157_6 ( .fault(fault), .net(N1157), .FEN(FEN[619]), .op(N1157_t6) );
fim FAN_N1157_7 ( .fault(fault), .net(N1157), .FEN(FEN[620]), .op(N1157_t7) );
fim FAN_N1157_8 ( .fault(fault), .net(N1157), .FEN(FEN[621]), .op(N1157_t8) );
fim FAN_N1157_9 ( .fault(fault), .net(N1157), .FEN(FEN[622]), .op(N1157_t9) );
fim FAN_N1173_0 ( .fault(fault), .net(N1173), .FEN(FEN[623]), .op(N1173_t0) );
fim FAN_N1173_1 ( .fault(fault), .net(N1173), .FEN(FEN[624]), .op(N1173_t1) );
fim FAN_N1173_2 ( .fault(fault), .net(N1173), .FEN(FEN[625]), .op(N1173_t2) );
fim FAN_N1173_3 ( .fault(fault), .net(N1173), .FEN(FEN[626]), .op(N1173_t3) );
fim FAN_N1178_0 ( .fault(fault), .net(N1178), .FEN(FEN[627]), .op(N1178_t0) );
fim FAN_N1178_1 ( .fault(fault), .net(N1178), .FEN(FEN[628]), .op(N1178_t1) );
fim FAN_N1178_2 ( .fault(fault), .net(N1178), .FEN(FEN[629]), .op(N1178_t2) );
fim FAN_N1178_3 ( .fault(fault), .net(N1178), .FEN(FEN[630]), .op(N1178_t3) );
fim FAN_N1178_4 ( .fault(fault), .net(N1178), .FEN(FEN[631]), .op(N1178_t4) );
fim FAN_N1200_0 ( .fault(fault), .net(N1200), .FEN(FEN[632]), .op(N1200_t0) );
fim FAN_N1200_1 ( .fault(fault), .net(N1200), .FEN(FEN[633]), .op(N1200_t1) );
fim FAN_N1200_2 ( .fault(fault), .net(N1200), .FEN(FEN[634]), .op(N1200_t2) );
fim FAN_N1200_3 ( .fault(fault), .net(N1200), .FEN(FEN[635]), .op(N1200_t3) );
fim FAN_N1205_0 ( .fault(fault), .net(N1205), .FEN(FEN[636]), .op(N1205_t0) );
fim FAN_N1205_1 ( .fault(fault), .net(N1205), .FEN(FEN[637]), .op(N1205_t1) );
fim FAN_N1205_2 ( .fault(fault), .net(N1205), .FEN(FEN[638]), .op(N1205_t2) );
fim FAN_N1205_3 ( .fault(fault), .net(N1205), .FEN(FEN[639]), .op(N1205_t3) );
fim FAN_N1251_0 ( .fault(fault), .net(N1251), .FEN(FEN[640]), .op(N1251_t0) );
fim FAN_N1251_1 ( .fault(fault), .net(N1251), .FEN(FEN[641]), .op(N1251_t1) );
fim FAN_N1254_0 ( .fault(fault), .net(N1254), .FEN(FEN[642]), .op(N1254_t0) );
fim FAN_N1254_1 ( .fault(fault), .net(N1254), .FEN(FEN[643]), .op(N1254_t1) );
fim FAN_N1257_0 ( .fault(fault), .net(N1257), .FEN(FEN[644]), .op(N1257_t0) );
fim FAN_N1257_1 ( .fault(fault), .net(N1257), .FEN(FEN[645]), .op(N1257_t1) );
fim FAN_N1260_0 ( .fault(fault), .net(N1260), .FEN(FEN[646]), .op(N1260_t0) );
fim FAN_N1260_1 ( .fault(fault), .net(N1260), .FEN(FEN[647]), .op(N1260_t1) );
fim FAN_N1263_0 ( .fault(fault), .net(N1263), .FEN(FEN[648]), .op(N1263_t0) );
fim FAN_N1263_1 ( .fault(fault), .net(N1263), .FEN(FEN[649]), .op(N1263_t1) );
fim FAN_N1266_0 ( .fault(fault), .net(N1266), .FEN(FEN[650]), .op(N1266_t0) );
fim FAN_N1266_1 ( .fault(fault), .net(N1266), .FEN(FEN[651]), .op(N1266_t1) );
fim FAN_N1216_0 ( .fault(fault), .net(N1216), .FEN(FEN[652]), .op(N1216_t0) );
fim FAN_N1216_1 ( .fault(fault), .net(N1216), .FEN(FEN[653]), .op(N1216_t1) );
fim FAN_N1591_0 ( .fault(fault), .net(N1591), .FEN(FEN[654]), .op(N1591_t0) );
fim FAN_N1591_1 ( .fault(fault), .net(N1591), .FEN(FEN[655]), .op(N1591_t1) );
fim FAN_N1591_2 ( .fault(fault), .net(N1591), .FEN(FEN[656]), .op(N1591_t2) );
fim FAN_N1591_3 ( .fault(fault), .net(N1591), .FEN(FEN[657]), .op(N1591_t3) );
fim FAN_N1502_0 ( .fault(fault), .net(N1502), .FEN(FEN[658]), .op(N1502_t0) );
fim FAN_N1502_1 ( .fault(fault), .net(N1502), .FEN(FEN[659]), .op(N1502_t1) );
fim FAN_N1502_2 ( .fault(fault), .net(N1502), .FEN(FEN[660]), .op(N1502_t2) );
fim FAN_N1506_0 ( .fault(fault), .net(N1506), .FEN(FEN[661]), .op(N1506_t0) );
fim FAN_N1506_1 ( .fault(fault), .net(N1506), .FEN(FEN[662]), .op(N1506_t1) );
fim FAN_N1506_2 ( .fault(fault), .net(N1506), .FEN(FEN[663]), .op(N1506_t2) );
fim FAN_N1513_0 ( .fault(fault), .net(N1513), .FEN(FEN[664]), .op(N1513_t0) );
fim FAN_N1513_1 ( .fault(fault), .net(N1513), .FEN(FEN[665]), .op(N1513_t1) );
fim FAN_N1516_0 ( .fault(fault), .net(N1516), .FEN(FEN[666]), .op(N1516_t0) );
fim FAN_N1516_1 ( .fault(fault), .net(N1516), .FEN(FEN[667]), .op(N1516_t1) );
fim FAN_N1510_0 ( .fault(fault), .net(N1510), .FEN(FEN[668]), .op(N1510_t0) );
fim FAN_N1510_1 ( .fault(fault), .net(N1510), .FEN(FEN[669]), .op(N1510_t1) );
fim FAN_N1499_0 ( .fault(fault), .net(N1499), .FEN(FEN[670]), .op(N1499_t0) );
fim FAN_N1499_1 ( .fault(fault), .net(N1499), .FEN(FEN[671]), .op(N1499_t1) );
fim FAN_N1496_0 ( .fault(fault), .net(N1496), .FEN(FEN[672]), .op(N1496_t0) );
fim FAN_N1496_1 ( .fault(fault), .net(N1496), .FEN(FEN[673]), .op(N1496_t1) );
fim FAN_N1553_0 ( .fault(fault), .net(N1553), .FEN(FEN[674]), .op(N1553_t0) );
fim FAN_N1553_1 ( .fault(fault), .net(N1553), .FEN(FEN[675]), .op(N1553_t1) );
fim FAN_N1553_2 ( .fault(fault), .net(N1553), .FEN(FEN[676]), .op(N1553_t2) );
fim FAN_N1557_0 ( .fault(fault), .net(N1557), .FEN(FEN[677]), .op(N1557_t0) );
fim FAN_N1557_1 ( .fault(fault), .net(N1557), .FEN(FEN[678]), .op(N1557_t1) );
fim FAN_N1557_2 ( .fault(fault), .net(N1557), .FEN(FEN[679]), .op(N1557_t2) );
fim FAN_N1561_0 ( .fault(fault), .net(N1561), .FEN(FEN[680]), .op(N1561_t0) );
fim FAN_N1561_1 ( .fault(fault), .net(N1561), .FEN(FEN[681]), .op(N1561_t1) );
fim FAN_N1588_0 ( .fault(fault), .net(N1588), .FEN(FEN[682]), .op(N1588_t0) );
fim FAN_N1588_1 ( .fault(fault), .net(N1588), .FEN(FEN[683]), .op(N1588_t1) );
fim FAN_N1578_0 ( .fault(fault), .net(N1578), .FEN(FEN[684]), .op(N1578_t0) );
fim FAN_N1578_1 ( .fault(fault), .net(N1578), .FEN(FEN[685]), .op(N1578_t1) );
fim FAN_N1582_0 ( .fault(fault), .net(N1582), .FEN(FEN[686]), .op(N1582_t0) );
fim FAN_N1582_1 ( .fault(fault), .net(N1582), .FEN(FEN[687]), .op(N1582_t1) );
fim FAN_N1585_0 ( .fault(fault), .net(N1585), .FEN(FEN[688]), .op(N1585_t0) );
fim FAN_N1585_1 ( .fault(fault), .net(N1585), .FEN(FEN[689]), .op(N1585_t1) );
fim FAN_N1596_0 ( .fault(fault), .net(N1596), .FEN(FEN[690]), .op(N1596_t0) );
fim FAN_N1596_1 ( .fault(fault), .net(N1596), .FEN(FEN[691]), .op(N1596_t1) );
fim FAN_N1596_2 ( .fault(fault), .net(N1596), .FEN(FEN[692]), .op(N1596_t2) );
fim FAN_N1606_0 ( .fault(fault), .net(N1606), .FEN(FEN[693]), .op(N1606_t0) );
fim FAN_N1606_1 ( .fault(fault), .net(N1606), .FEN(FEN[694]), .op(N1606_t1) );
fim FAN_N1606_2 ( .fault(fault), .net(N1606), .FEN(FEN[695]), .op(N1606_t2) );
fim FAN_N1606_3 ( .fault(fault), .net(N1606), .FEN(FEN[696]), .op(N1606_t3) );
fim FAN_N1606_4 ( .fault(fault), .net(N1606), .FEN(FEN[697]), .op(N1606_t4) );
fim FAN_N1600_0 ( .fault(fault), .net(N1600), .FEN(FEN[698]), .op(N1600_t0) );
fim FAN_N1600_1 ( .fault(fault), .net(N1600), .FEN(FEN[699]), .op(N1600_t1) );
fim FAN_N1600_2 ( .fault(fault), .net(N1600), .FEN(FEN[700]), .op(N1600_t2) );
fim FAN_N1600_3 ( .fault(fault), .net(N1600), .FEN(FEN[701]), .op(N1600_t3) );
fim FAN_N1600_4 ( .fault(fault), .net(N1600), .FEN(FEN[702]), .op(N1600_t4) );
fim FAN_N1642_0 ( .fault(fault), .net(N1642), .FEN(FEN[703]), .op(N1642_t0) );
fim FAN_N1642_1 ( .fault(fault), .net(N1642), .FEN(FEN[704]), .op(N1642_t1) );
fim FAN_N1642_2 ( .fault(fault), .net(N1642), .FEN(FEN[705]), .op(N1642_t2) );
fim FAN_N1642_3 ( .fault(fault), .net(N1642), .FEN(FEN[706]), .op(N1642_t3) );
fim FAN_N1647_0 ( .fault(fault), .net(N1647), .FEN(FEN[707]), .op(N1647_t0) );
fim FAN_N1647_1 ( .fault(fault), .net(N1647), .FEN(FEN[708]), .op(N1647_t1) );
fim FAN_N1647_2 ( .fault(fault), .net(N1647), .FEN(FEN[709]), .op(N1647_t2) );
fim FAN_N1637_0 ( .fault(fault), .net(N1637), .FEN(FEN[710]), .op(N1637_t0) );
fim FAN_N1637_1 ( .fault(fault), .net(N1637), .FEN(FEN[711]), .op(N1637_t1) );
fim FAN_N1637_2 ( .fault(fault), .net(N1637), .FEN(FEN[712]), .op(N1637_t2) );
fim FAN_N1637_3 ( .fault(fault), .net(N1637), .FEN(FEN[713]), .op(N1637_t3) );
fim FAN_N1624_0 ( .fault(fault), .net(N1624), .FEN(FEN[714]), .op(N1624_t0) );
fim FAN_N1624_1 ( .fault(fault), .net(N1624), .FEN(FEN[715]), .op(N1624_t1) );
fim FAN_N1624_2 ( .fault(fault), .net(N1624), .FEN(FEN[716]), .op(N1624_t2) );
fim FAN_N1619_0 ( .fault(fault), .net(N1619), .FEN(FEN[717]), .op(N1619_t0) );
fim FAN_N1619_1 ( .fault(fault), .net(N1619), .FEN(FEN[718]), .op(N1619_t1) );
fim FAN_N1619_2 ( .fault(fault), .net(N1619), .FEN(FEN[719]), .op(N1619_t2) );
fim FAN_N1619_3 ( .fault(fault), .net(N1619), .FEN(FEN[720]), .op(N1619_t3) );
fim FAN_N1615_0 ( .fault(fault), .net(N1615), .FEN(FEN[721]), .op(N1615_t0) );
fim FAN_N1615_1 ( .fault(fault), .net(N1615), .FEN(FEN[722]), .op(N1615_t1) );
fim FAN_N1615_2 ( .fault(fault), .net(N1615), .FEN(FEN[723]), .op(N1615_t2) );
fim FAN_N496_0 ( .fault(fault), .net(N496), .FEN(FEN[724]), .op(N496_t0) );
fim FAN_N496_1 ( .fault(fault), .net(N496), .FEN(FEN[725]), .op(N496_t1) );
fim FAN_N224_0 ( .fault(fault), .net(N224), .FEN(FEN[726]), .op(N224_t0) );
fim FAN_N224_1 ( .fault(fault), .net(N224), .FEN(FEN[727]), .op(N224_t1) );
fim FAN_N1612_0 ( .fault(fault), .net(N1612), .FEN(FEN[728]), .op(N1612_t0) );
fim FAN_N1612_1 ( .fault(fault), .net(N1612), .FEN(FEN[729]), .op(N1612_t1) );
fim FAN_N1628_0 ( .fault(fault), .net(N1628), .FEN(FEN[730]), .op(N1628_t0) );
fim FAN_N1628_1 ( .fault(fault), .net(N1628), .FEN(FEN[731]), .op(N1628_t1) );
fim FAN_N1631_0 ( .fault(fault), .net(N1631), .FEN(FEN[732]), .op(N1631_t0) );
fim FAN_N1631_1 ( .fault(fault), .net(N1631), .FEN(FEN[733]), .op(N1631_t1) );
fim FAN_N1634_0 ( .fault(fault), .net(N1634), .FEN(FEN[734]), .op(N1634_t0) );
fim FAN_N1634_1 ( .fault(fault), .net(N1634), .FEN(FEN[735]), .op(N1634_t1) );
fim FAN_N727_0 ( .fault(fault), .net(N727), .FEN(FEN[736]), .op(N727_t0) );
fim FAN_N727_1 ( .fault(fault), .net(N727), .FEN(FEN[737]), .op(N727_t1) );
fim FAN_N1651_0 ( .fault(fault), .net(N1651), .FEN(FEN[738]), .op(N1651_t0) );
fim FAN_N1651_1 ( .fault(fault), .net(N1651), .FEN(FEN[739]), .op(N1651_t1) );
fim FAN_N1651_2 ( .fault(fault), .net(N1651), .FEN(FEN[740]), .op(N1651_t2) );
fim FAN_N1651_3 ( .fault(fault), .net(N1651), .FEN(FEN[741]), .op(N1651_t3) );
fim FAN_N730_0 ( .fault(fault), .net(N730), .FEN(FEN[742]), .op(N730_t0) );
fim FAN_N730_1 ( .fault(fault), .net(N730), .FEN(FEN[743]), .op(N730_t1) );
fim FAN_N1656_0 ( .fault(fault), .net(N1656), .FEN(FEN[744]), .op(N1656_t0) );
fim FAN_N1656_1 ( .fault(fault), .net(N1656), .FEN(FEN[745]), .op(N1656_t1) );
fim FAN_N1656_2 ( .fault(fault), .net(N1656), .FEN(FEN[746]), .op(N1656_t2) );
fim FAN_N1686_0 ( .fault(fault), .net(N1686), .FEN(FEN[747]), .op(N1686_t0) );
fim FAN_N1686_1 ( .fault(fault), .net(N1686), .FEN(FEN[748]), .op(N1686_t1) );
fim FAN_N1686_2 ( .fault(fault), .net(N1686), .FEN(FEN[749]), .op(N1686_t2) );
fim FAN_N1708_0 ( .fault(fault), .net(N1708), .FEN(FEN[750]), .op(N1708_t0) );
fim FAN_N1708_1 ( .fault(fault), .net(N1708), .FEN(FEN[751]), .op(N1708_t1) );
fim FAN_N1676_0 ( .fault(fault), .net(N1676), .FEN(FEN[752]), .op(N1676_t0) );
fim FAN_N1676_1 ( .fault(fault), .net(N1676), .FEN(FEN[753]), .op(N1676_t1) );
fim FAN_N1676_2 ( .fault(fault), .net(N1676), .FEN(FEN[754]), .op(N1676_t2) );
fim FAN_N1676_3 ( .fault(fault), .net(N1676), .FEN(FEN[755]), .op(N1676_t3) );
fim FAN_N1681_0 ( .fault(fault), .net(N1681), .FEN(FEN[756]), .op(N1681_t0) );
fim FAN_N1681_1 ( .fault(fault), .net(N1681), .FEN(FEN[757]), .op(N1681_t1) );
fim FAN_N1681_2 ( .fault(fault), .net(N1681), .FEN(FEN[758]), .op(N1681_t2) );
fim FAN_N1681_3 ( .fault(fault), .net(N1681), .FEN(FEN[759]), .op(N1681_t3) );
fim FAN_N1690_0 ( .fault(fault), .net(N1690), .FEN(FEN[760]), .op(N1690_t0) );
fim FAN_N1690_1 ( .fault(fault), .net(N1690), .FEN(FEN[761]), .op(N1690_t1) );
fim FAN_N533_0 ( .fault(fault), .net(N533), .FEN(FEN[762]), .op(N533_t0) );
fim FAN_N533_1 ( .fault(fault), .net(N533), .FEN(FEN[763]), .op(N533_t1) );
fim FAN_N533_2 ( .fault(fault), .net(N533), .FEN(FEN[764]), .op(N533_t2) );
fim FAN_N1848_0 ( .fault(fault), .net(N1848), .FEN(FEN[765]), .op(N1848_t0) );
fim FAN_N1848_1 ( .fault(fault), .net(N1848), .FEN(FEN[766]), .op(N1848_t1) );
fim FAN_N1848_2 ( .fault(fault), .net(N1848), .FEN(FEN[767]), .op(N1848_t2) );
fim FAN_N1852_0 ( .fault(fault), .net(N1852), .FEN(FEN[768]), .op(N1852_t0) );
fim FAN_N1852_1 ( .fault(fault), .net(N1852), .FEN(FEN[769]), .op(N1852_t1) );
fim FAN_N1852_2 ( .fault(fault), .net(N1852), .FEN(FEN[770]), .op(N1852_t2) );
fim FAN_N1856_0 ( .fault(fault), .net(N1856), .FEN(FEN[771]), .op(N1856_t0) );
fim FAN_N1856_1 ( .fault(fault), .net(N1856), .FEN(FEN[772]), .op(N1856_t1) );
fim FAN_N1856_2 ( .fault(fault), .net(N1856), .FEN(FEN[773]), .op(N1856_t2) );
fim FAN_N1856_3 ( .fault(fault), .net(N1856), .FEN(FEN[774]), .op(N1856_t3) );
fim FAN_N1856_4 ( .fault(fault), .net(N1856), .FEN(FEN[775]), .op(N1856_t4) );
fim FAN_N1856_5 ( .fault(fault), .net(N1856), .FEN(FEN[776]), .op(N1856_t5) );
fim FAN_N1863_0 ( .fault(fault), .net(N1863), .FEN(FEN[777]), .op(N1863_t0) );
fim FAN_N1863_1 ( .fault(fault), .net(N1863), .FEN(FEN[778]), .op(N1863_t1) );
fim FAN_N1863_2 ( .fault(fault), .net(N1863), .FEN(FEN[779]), .op(N1863_t2) );
fim FAN_N1863_3 ( .fault(fault), .net(N1863), .FEN(FEN[780]), .op(N1863_t3) );
fim FAN_N1863_4 ( .fault(fault), .net(N1863), .FEN(FEN[781]), .op(N1863_t4) );
fim FAN_N1863_5 ( .fault(fault), .net(N1863), .FEN(FEN[782]), .op(N1863_t5) );
fim FAN_N1870_0 ( .fault(fault), .net(N1870), .FEN(FEN[783]), .op(N1870_t0) );
fim FAN_N1870_1 ( .fault(fault), .net(N1870), .FEN(FEN[784]), .op(N1870_t1) );
fim FAN_N1870_2 ( .fault(fault), .net(N1870), .FEN(FEN[785]), .op(N1870_t2) );
fim FAN_N1870_3 ( .fault(fault), .net(N1870), .FEN(FEN[786]), .op(N1870_t3) );
fim FAN_N1875_0 ( .fault(fault), .net(N1875), .FEN(FEN[787]), .op(N1875_t0) );
fim FAN_N1875_1 ( .fault(fault), .net(N1875), .FEN(FEN[788]), .op(N1875_t1) );
fim FAN_N1875_2 ( .fault(fault), .net(N1875), .FEN(FEN[789]), .op(N1875_t2) );
fim FAN_N1875_3 ( .fault(fault), .net(N1875), .FEN(FEN[790]), .op(N1875_t3) );
fim FAN_N1880_0 ( .fault(fault), .net(N1880), .FEN(FEN[791]), .op(N1880_t0) );
fim FAN_N1880_1 ( .fault(fault), .net(N1880), .FEN(FEN[792]), .op(N1880_t1) );
fim FAN_N1880_2 ( .fault(fault), .net(N1880), .FEN(FEN[793]), .op(N1880_t2) );
fim FAN_N1880_3 ( .fault(fault), .net(N1880), .FEN(FEN[794]), .op(N1880_t3) );
fim FAN_N1778_0 ( .fault(fault), .net(N1778), .FEN(FEN[795]), .op(N1778_t0) );
fim FAN_N1778_1 ( .fault(fault), .net(N1778), .FEN(FEN[796]), .op(N1778_t1) );
fim FAN_N1781_0 ( .fault(fault), .net(N1781), .FEN(FEN[797]), .op(N1781_t0) );
fim FAN_N1781_1 ( .fault(fault), .net(N1781), .FEN(FEN[798]), .op(N1781_t1) );
fim FAN_N1773_0 ( .fault(fault), .net(N1773), .FEN(FEN[799]), .op(N1773_t0) );
fim FAN_N1773_1 ( .fault(fault), .net(N1773), .FEN(FEN[800]), .op(N1773_t1) );
fim FAN_N1770_0 ( .fault(fault), .net(N1770), .FEN(FEN[801]), .op(N1770_t0) );
fim FAN_N1770_1 ( .fault(fault), .net(N1770), .FEN(FEN[802]), .op(N1770_t1) );
fim FAN_N1801_0 ( .fault(fault), .net(N1801), .FEN(FEN[803]), .op(N1801_t0) );
fim FAN_N1801_1 ( .fault(fault), .net(N1801), .FEN(FEN[804]), .op(N1801_t1) );
fim FAN_N1804_0 ( .fault(fault), .net(N1804), .FEN(FEN[805]), .op(N1804_t0) );
fim FAN_N1804_1 ( .fault(fault), .net(N1804), .FEN(FEN[806]), .op(N1804_t1) );
fim FAN_N1798_0 ( .fault(fault), .net(N1798), .FEN(FEN[807]), .op(N1798_t0) );
fim FAN_N1798_1 ( .fault(fault), .net(N1798), .FEN(FEN[808]), .op(N1798_t1) );
fim FAN_N1795_0 ( .fault(fault), .net(N1795), .FEN(FEN[809]), .op(N1795_t0) );
fim FAN_N1795_1 ( .fault(fault), .net(N1795), .FEN(FEN[810]), .op(N1795_t1) );
fim FAN_N1897_0 ( .fault(fault), .net(N1897), .FEN(FEN[811]), .op(N1897_t0) );
fim FAN_N1897_1 ( .fault(fault), .net(N1897), .FEN(FEN[812]), .op(N1897_t1) );
fim FAN_N1894_0 ( .fault(fault), .net(N1894), .FEN(FEN[813]), .op(N1894_t0) );
fim FAN_N1894_1 ( .fault(fault), .net(N1894), .FEN(FEN[814]), .op(N1894_t1) );
fim FAN_N40_0 ( .fault(fault), .net(N40), .FEN(FEN[815]), .op(N40_t0) );
fim FAN_N40_1 ( .fault(fault), .net(N40), .FEN(FEN[816]), .op(N40_t1) );
fim FAN_N1827_0 ( .fault(fault), .net(N1827), .FEN(FEN[817]), .op(N1827_t0) );
fim FAN_N1827_1 ( .fault(fault), .net(N1827), .FEN(FEN[818]), .op(N1827_t1) );
fim FAN_N1824_0 ( .fault(fault), .net(N1824), .FEN(FEN[819]), .op(N1824_t0) );
fim FAN_N1824_1 ( .fault(fault), .net(N1824), .FEN(FEN[820]), .op(N1824_t1) );
fim FAN_N1885_0 ( .fault(fault), .net(N1885), .FEN(FEN[821]), .op(N1885_t0) );
fim FAN_N1885_1 ( .fault(fault), .net(N1885), .FEN(FEN[822]), .op(N1885_t1) );
fim FAN_N1888_0 ( .fault(fault), .net(N1888), .FEN(FEN[823]), .op(N1888_t0) );
fim FAN_N1888_1 ( .fault(fault), .net(N1888), .FEN(FEN[824]), .op(N1888_t1) );
fim FAN_N1942_0 ( .fault(fault), .net(N1942), .FEN(FEN[825]), .op(N1942_t0) );
fim FAN_N1942_1 ( .fault(fault), .net(N1942), .FEN(FEN[826]), .op(N1942_t1) );
fim FAN_N1945_0 ( .fault(fault), .net(N1945), .FEN(FEN[827]), .op(N1945_t0) );
fim FAN_N1945_1 ( .fault(fault), .net(N1945), .FEN(FEN[828]), .op(N1945_t1) );
fim FAN_N1948_0 ( .fault(fault), .net(N1948), .FEN(FEN[829]), .op(N1948_t0) );
fim FAN_N1948_1 ( .fault(fault), .net(N1948), .FEN(FEN[830]), .op(N1948_t1) );
fim FAN_N1951_0 ( .fault(fault), .net(N1951), .FEN(FEN[831]), .op(N1951_t0) );
fim FAN_N1951_1 ( .fault(fault), .net(N1951), .FEN(FEN[832]), .op(N1951_t1) );
fim FAN_N1954_0 ( .fault(fault), .net(N1954), .FEN(FEN[833]), .op(N1954_t0) );
fim FAN_N1954_1 ( .fault(fault), .net(N1954), .FEN(FEN[834]), .op(N1954_t1) );
fim FAN_N1836_0 ( .fault(fault), .net(N1836), .FEN(FEN[835]), .op(N1836_t0) );
fim FAN_N1836_1 ( .fault(fault), .net(N1836), .FEN(FEN[836]), .op(N1836_t1) );
fim FAN_N1836_2 ( .fault(fault), .net(N1836), .FEN(FEN[837]), .op(N1836_t2) );
fim FAN_N1836_3 ( .fault(fault), .net(N1836), .FEN(FEN[838]), .op(N1836_t3) );
fim FAN_N1833_0 ( .fault(fault), .net(N1833), .FEN(FEN[839]), .op(N1833_t0) );
fim FAN_N1833_1 ( .fault(fault), .net(N1833), .FEN(FEN[840]), .op(N1833_t1) );
fim FAN_N1841_0 ( .fault(fault), .net(N1841), .FEN(FEN[841]), .op(N1841_t0) );
fim FAN_N1841_1 ( .fault(fault), .net(N1841), .FEN(FEN[842]), .op(N1841_t1) );
fim FAN_N1841_2 ( .fault(fault), .net(N1841), .FEN(FEN[843]), .op(N1841_t2) );
fim FAN_N1841_3 ( .fault(fault), .net(N1841), .FEN(FEN[844]), .op(N1841_t3) );
fim FAN_N1841_4 ( .fault(fault), .net(N1841), .FEN(FEN[845]), .op(N1841_t4) );
fim FAN_N1841_5 ( .fault(fault), .net(N1841), .FEN(FEN[846]), .op(N1841_t5) );
fim FAN_N1936_0 ( .fault(fault), .net(N1936), .FEN(FEN[847]), .op(N1936_t0) );
fim FAN_N1936_1 ( .fault(fault), .net(N1936), .FEN(FEN[848]), .op(N1936_t1) );
fim FAN_N1957_0 ( .fault(fault), .net(N1957), .FEN(FEN[849]), .op(N1957_t0) );
fim FAN_N1957_1 ( .fault(fault), .net(N1957), .FEN(FEN[850]), .op(N1957_t1) );
fim FAN_N1960_0 ( .fault(fault), .net(N1960), .FEN(FEN[851]), .op(N1960_t0) );
fim FAN_N1960_1 ( .fault(fault), .net(N1960), .FEN(FEN[852]), .op(N1960_t1) );
fim FAN_N1963_0 ( .fault(fault), .net(N1963), .FEN(FEN[853]), .op(N1963_t0) );
fim FAN_N1963_1 ( .fault(fault), .net(N1963), .FEN(FEN[854]), .op(N1963_t1) );
fim FAN_N1966_0 ( .fault(fault), .net(N1966), .FEN(FEN[855]), .op(N1966_t0) );
fim FAN_N1966_1 ( .fault(fault), .net(N1966), .FEN(FEN[856]), .op(N1966_t1) );
fim FAN_N2046_0 ( .fault(fault), .net(N2046), .FEN(FEN[857]), .op(N2046_t0) );
fim FAN_N2046_1 ( .fault(fault), .net(N2046), .FEN(FEN[858]), .op(N2046_t1) );
fim FAN_N2049_0 ( .fault(fault), .net(N2049), .FEN(FEN[859]), .op(N2049_t0) );
fim FAN_N2049_1 ( .fault(fault), .net(N2049), .FEN(FEN[860]), .op(N2049_t1) );
fim FAN_N2052_0 ( .fault(fault), .net(N2052), .FEN(FEN[861]), .op(N2052_t0) );
fim FAN_N2052_1 ( .fault(fault), .net(N2052), .FEN(FEN[862]), .op(N2052_t1) );
fim FAN_N2055_0 ( .fault(fault), .net(N2055), .FEN(FEN[863]), .op(N2055_t0) );
fim FAN_N2055_1 ( .fault(fault), .net(N2055), .FEN(FEN[864]), .op(N2055_t1) );
fim FAN_N2058_0 ( .fault(fault), .net(N2058), .FEN(FEN[865]), .op(N2058_t0) );
fim FAN_N2058_1 ( .fault(fault), .net(N2058), .FEN(FEN[866]), .op(N2058_t1) );
fim FAN_N2061_0 ( .fault(fault), .net(N2061), .FEN(FEN[867]), .op(N2061_t0) );
fim FAN_N2061_1 ( .fault(fault), .net(N2061), .FEN(FEN[868]), .op(N2061_t1) );
fim FAN_N2064_0 ( .fault(fault), .net(N2064), .FEN(FEN[869]), .op(N2064_t0) );
fim FAN_N2064_1 ( .fault(fault), .net(N2064), .FEN(FEN[870]), .op(N2064_t1) );
fim FAN_N2067_0 ( .fault(fault), .net(N2067), .FEN(FEN[871]), .op(N2067_t0) );
fim FAN_N2067_1 ( .fault(fault), .net(N2067), .FEN(FEN[872]), .op(N2067_t1) );
fim FAN_N2070_0 ( .fault(fault), .net(N2070), .FEN(FEN[873]), .op(N2070_t0) );
fim FAN_N2070_1 ( .fault(fault), .net(N2070), .FEN(FEN[874]), .op(N2070_t1) );
fim FAN_N2073_0 ( .fault(fault), .net(N2073), .FEN(FEN[875]), .op(N2073_t0) );
fim FAN_N2073_1 ( .fault(fault), .net(N2073), .FEN(FEN[876]), .op(N2073_t1) );
fim FAN_N2076_0 ( .fault(fault), .net(N2076), .FEN(FEN[877]), .op(N2076_t0) );
fim FAN_N2076_1 ( .fault(fault), .net(N2076), .FEN(FEN[878]), .op(N2076_t1) );
fim FAN_N2079_0 ( .fault(fault), .net(N2079), .FEN(FEN[879]), .op(N2079_t0) );
fim FAN_N2079_1 ( .fault(fault), .net(N2079), .FEN(FEN[880]), .op(N2079_t1) );
fim FAN_N2095_0 ( .fault(fault), .net(N2095), .FEN(FEN[881]), .op(N2095_t0) );
fim FAN_N2095_1 ( .fault(fault), .net(N2095), .FEN(FEN[882]), .op(N2095_t1) );
fim FAN_N2098_0 ( .fault(fault), .net(N2098), .FEN(FEN[883]), .op(N2098_t0) );
fim FAN_N2098_1 ( .fault(fault), .net(N2098), .FEN(FEN[884]), .op(N2098_t1) );
fim FAN_N2101_0 ( .fault(fault), .net(N2101), .FEN(FEN[885]), .op(N2101_t0) );
fim FAN_N2101_1 ( .fault(fault), .net(N2101), .FEN(FEN[886]), .op(N2101_t1) );
fim FAN_N2104_0 ( .fault(fault), .net(N2104), .FEN(FEN[887]), .op(N2104_t0) );
fim FAN_N2104_1 ( .fault(fault), .net(N2104), .FEN(FEN[888]), .op(N2104_t1) );
fim FAN_N2107_0 ( .fault(fault), .net(N2107), .FEN(FEN[889]), .op(N2107_t0) );
fim FAN_N2107_1 ( .fault(fault), .net(N2107), .FEN(FEN[890]), .op(N2107_t1) );
fim FAN_N2110_0 ( .fault(fault), .net(N2110), .FEN(FEN[891]), .op(N2110_t0) );
fim FAN_N2110_1 ( .fault(fault), .net(N2110), .FEN(FEN[892]), .op(N2110_t1) );
fim FAN_N2120_0 ( .fault(fault), .net(N2120), .FEN(FEN[893]), .op(N2120_t0) );
fim FAN_N2120_1 ( .fault(fault), .net(N2120), .FEN(FEN[894]), .op(N2120_t1) );
fim FAN_N2120_2 ( .fault(fault), .net(N2120), .FEN(FEN[895]), .op(N2120_t2) );
fim FAN_N2120_3 ( .fault(fault), .net(N2120), .FEN(FEN[896]), .op(N2120_t3) );
fim FAN_N2113_0 ( .fault(fault), .net(N2113), .FEN(FEN[897]), .op(N2113_t0) );
fim FAN_N2113_1 ( .fault(fault), .net(N2113), .FEN(FEN[898]), .op(N2113_t1) );
fim FAN_N2113_2 ( .fault(fault), .net(N2113), .FEN(FEN[899]), .op(N2113_t2) );
fim FAN_N2113_3 ( .fault(fault), .net(N2113), .FEN(FEN[900]), .op(N2113_t3) );
fim FAN_N2113_4 ( .fault(fault), .net(N2113), .FEN(FEN[901]), .op(N2113_t4) );
fim FAN_N2185_0 ( .fault(fault), .net(N2185), .FEN(FEN[902]), .op(N2185_t0) );
fim FAN_N2185_1 ( .fault(fault), .net(N2185), .FEN(FEN[903]), .op(N2185_t1) );
fim FAN_N2188_0 ( .fault(fault), .net(N2188), .FEN(FEN[904]), .op(N2188_t0) );
fim FAN_N2188_1 ( .fault(fault), .net(N2188), .FEN(FEN[905]), .op(N2188_t1) );
fim FAN_N2191_0 ( .fault(fault), .net(N2191), .FEN(FEN[906]), .op(N2191_t0) );
fim FAN_N2191_1 ( .fault(fault), .net(N2191), .FEN(FEN[907]), .op(N2191_t1) );
fim FAN_N2194_0 ( .fault(fault), .net(N2194), .FEN(FEN[908]), .op(N2194_t0) );
fim FAN_N2194_1 ( .fault(fault), .net(N2194), .FEN(FEN[909]), .op(N2194_t1) );
fim FAN_N2201_0 ( .fault(fault), .net(N2201), .FEN(FEN[910]), .op(N2201_t0) );
fim FAN_N2201_1 ( .fault(fault), .net(N2201), .FEN(FEN[911]), .op(N2201_t1) );
fim FAN_N2204_0 ( .fault(fault), .net(N2204), .FEN(FEN[912]), .op(N2204_t0) );
fim FAN_N2204_1 ( .fault(fault), .net(N2204), .FEN(FEN[913]), .op(N2204_t1) );
fim FAN_N2207_0 ( .fault(fault), .net(N2207), .FEN(FEN[914]), .op(N2207_t0) );
fim FAN_N2207_1 ( .fault(fault), .net(N2207), .FEN(FEN[915]), .op(N2207_t1) );
fim FAN_N2210_0 ( .fault(fault), .net(N2210), .FEN(FEN[916]), .op(N2210_t0) );
fim FAN_N2210_1 ( .fault(fault), .net(N2210), .FEN(FEN[917]), .op(N2210_t1) );
fim FAN_N2213_0 ( .fault(fault), .net(N2213), .FEN(FEN[918]), .op(N2213_t0) );
fim FAN_N2213_1 ( .fault(fault), .net(N2213), .FEN(FEN[919]), .op(N2213_t1) );
fim FAN_N2266_0 ( .fault(fault), .net(N2266), .FEN(FEN[920]), .op(N2266_t0) );
fim FAN_N2266_1 ( .fault(fault), .net(N2266), .FEN(FEN[921]), .op(N2266_t1) );
fim FAN_N2269_0 ( .fault(fault), .net(N2269), .FEN(FEN[922]), .op(N2269_t0) );
fim FAN_N2269_1 ( .fault(fault), .net(N2269), .FEN(FEN[923]), .op(N2269_t1) );
fim FAN_N2219_0 ( .fault(fault), .net(N2219), .FEN(FEN[924]), .op(N2219_t0) );
fim FAN_N2219_1 ( .fault(fault), .net(N2219), .FEN(FEN[925]), .op(N2219_t1) );
fim FAN_N2216_0 ( .fault(fault), .net(N2216), .FEN(FEN[926]), .op(N2216_t0) );
fim FAN_N2216_1 ( .fault(fault), .net(N2216), .FEN(FEN[927]), .op(N2216_t1) );
fim FAN_N2128_0 ( .fault(fault), .net(N2128), .FEN(FEN[928]), .op(N2128_t0) );
fim FAN_N2128_1 ( .fault(fault), .net(N2128), .FEN(FEN[929]), .op(N2128_t1) );
fim FAN_N2128_2 ( .fault(fault), .net(N2128), .FEN(FEN[930]), .op(N2128_t2) );
fim FAN_N2128_3 ( .fault(fault), .net(N2128), .FEN(FEN[931]), .op(N2128_t3) );
fim FAN_N2128_4 ( .fault(fault), .net(N2128), .FEN(FEN[932]), .op(N2128_t4) );
fim FAN_N2128_5 ( .fault(fault), .net(N2128), .FEN(FEN[933]), .op(N2128_t5) );
fim FAN_N2135_0 ( .fault(fault), .net(N2135), .FEN(FEN[934]), .op(N2135_t0) );
fim FAN_N2135_1 ( .fault(fault), .net(N2135), .FEN(FEN[935]), .op(N2135_t1) );
fim FAN_N2135_2 ( .fault(fault), .net(N2135), .FEN(FEN[936]), .op(N2135_t2) );
fim FAN_N2135_3 ( .fault(fault), .net(N2135), .FEN(FEN[937]), .op(N2135_t3) );
fim FAN_N2135_4 ( .fault(fault), .net(N2135), .FEN(FEN[938]), .op(N2135_t4) );
fim FAN_N2144_0 ( .fault(fault), .net(N2144), .FEN(FEN[939]), .op(N2144_t0) );
fim FAN_N2144_1 ( .fault(fault), .net(N2144), .FEN(FEN[940]), .op(N2144_t1) );
fim FAN_N2141_0 ( .fault(fault), .net(N2141), .FEN(FEN[941]), .op(N2141_t0) );
fim FAN_N2141_1 ( .fault(fault), .net(N2141), .FEN(FEN[942]), .op(N2141_t1) );
fim FAN_N2150_0 ( .fault(fault), .net(N2150), .FEN(FEN[943]), .op(N2150_t0) );
fim FAN_N2150_1 ( .fault(fault), .net(N2150), .FEN(FEN[944]), .op(N2150_t1) );
fim FAN_N2147_0 ( .fault(fault), .net(N2147), .FEN(FEN[945]), .op(N2147_t0) );
fim FAN_N2147_1 ( .fault(fault), .net(N2147), .FEN(FEN[946]), .op(N2147_t1) );
fim FAN_N2197_0 ( .fault(fault), .net(N2197), .FEN(FEN[947]), .op(N2197_t0) );
fim FAN_N2197_1 ( .fault(fault), .net(N2197), .FEN(FEN[948]), .op(N2197_t1) );
fim FAN_N2291_0 ( .fault(fault), .net(N2291), .FEN(FEN[949]), .op(N2291_t0) );
fim FAN_N2291_1 ( .fault(fault), .net(N2291), .FEN(FEN[950]), .op(N2291_t1) );
fim FAN_N2294_0 ( .fault(fault), .net(N2294), .FEN(FEN[951]), .op(N2294_t0) );
fim FAN_N2294_1 ( .fault(fault), .net(N2294), .FEN(FEN[952]), .op(N2294_t1) );
fim FAN_N2250_0 ( .fault(fault), .net(N2250), .FEN(FEN[953]), .op(N2250_t0) );
fim FAN_N2250_1 ( .fault(fault), .net(N2250), .FEN(FEN[954]), .op(N2250_t1) );
fim FAN_N2359_0 ( .fault(fault), .net(N2359), .FEN(FEN[955]), .op(N2359_t0) );
fim FAN_N2359_1 ( .fault(fault), .net(N2359), .FEN(FEN[956]), .op(N2359_t1) );
fim FAN_N2377_0 ( .fault(fault), .net(N2377), .FEN(FEN[957]), .op(N2377_t0) );
fim FAN_N2377_1 ( .fault(fault), .net(N2377), .FEN(FEN[958]), .op(N2377_t1) );
fim FAN_N2377_2 ( .fault(fault), .net(N2377), .FEN(FEN[959]), .op(N2377_t2) );
fim FAN_N2377_3 ( .fault(fault), .net(N2377), .FEN(FEN[960]), .op(N2377_t3) );
fim FAN_N1891_0 ( .fault(fault), .net(N1891), .FEN(FEN[961]), .op(N1891_t0) );
fim FAN_N1891_1 ( .fault(fault), .net(N1891), .FEN(FEN[962]), .op(N1891_t1) );
fim FAN_N2382_0 ( .fault(fault), .net(N2382), .FEN(FEN[963]), .op(N2382_t0) );
fim FAN_N2382_1 ( .fault(fault), .net(N2382), .FEN(FEN[964]), .op(N2382_t1) );
fim FAN_N2382_2 ( .fault(fault), .net(N2382), .FEN(FEN[965]), .op(N2382_t2) );
fim FAN_N2434_0 ( .fault(fault), .net(N2434), .FEN(FEN[966]), .op(N2434_t0) );
fim FAN_N2434_1 ( .fault(fault), .net(N2434), .FEN(FEN[967]), .op(N2434_t1) );
fim FAN_N2437_0 ( .fault(fault), .net(N2437), .FEN(FEN[968]), .op(N2437_t0) );
fim FAN_N2437_1 ( .fault(fault), .net(N2437), .FEN(FEN[969]), .op(N2437_t1) );
fim FAN_N2368_0 ( .fault(fault), .net(N2368), .FEN(FEN[970]), .op(N2368_t0) );
fim FAN_N2368_1 ( .fault(fault), .net(N2368), .FEN(FEN[971]), .op(N2368_t1) );
fim FAN_N2368_2 ( .fault(fault), .net(N2368), .FEN(FEN[972]), .op(N2368_t2) );
fim FAN_N2454_0 ( .fault(fault), .net(N2454), .FEN(FEN[973]), .op(N2454_t0) );
fim FAN_N2454_1 ( .fault(fault), .net(N2454), .FEN(FEN[974]), .op(N2454_t1) );
fim FAN_N2472_0 ( .fault(fault), .net(N2472), .FEN(FEN[975]), .op(N2472_t0) );
fim FAN_N2472_1 ( .fault(fault), .net(N2472), .FEN(FEN[976]), .op(N2472_t1) );
fim FAN_N2391_0 ( .fault(fault), .net(N2391), .FEN(FEN[977]), .op(N2391_t0) );
fim FAN_N2391_1 ( .fault(fault), .net(N2391), .FEN(FEN[978]), .op(N2391_t1) );
fim FAN_N2391_2 ( .fault(fault), .net(N2391), .FEN(FEN[979]), .op(N2391_t2) );
fim FAN_N2395_0 ( .fault(fault), .net(N2395), .FEN(FEN[980]), .op(N2395_t0) );
fim FAN_N2395_1 ( .fault(fault), .net(N2395), .FEN(FEN[981]), .op(N2395_t1) );
fim FAN_N2395_2 ( .fault(fault), .net(N2395), .FEN(FEN[982]), .op(N2395_t2) );
fim FAN_N2395_3 ( .fault(fault), .net(N2395), .FEN(FEN[983]), .op(N2395_t3) );
fim FAN_N2521_0 ( .fault(fault), .net(N2521), .FEN(FEN[984]), .op(N2521_t0) );
fim FAN_N2521_1 ( .fault(fault), .net(N2521), .FEN(FEN[985]), .op(N2521_t1) );
fim FAN_N2475_0 ( .fault(fault), .net(N2475), .FEN(FEN[986]), .op(N2475_t0) );
fim FAN_N2475_1 ( .fault(fault), .net(N2475), .FEN(FEN[987]), .op(N2475_t1) );
fim FAN_N2478_0 ( .fault(fault), .net(N2478), .FEN(FEN[988]), .op(N2478_t0) );
fim FAN_N2478_1 ( .fault(fault), .net(N2478), .FEN(FEN[989]), .op(N2478_t1) );
fim FAN_N2481_0 ( .fault(fault), .net(N2481), .FEN(FEN[990]), .op(N2481_t0) );
fim FAN_N2481_1 ( .fault(fault), .net(N2481), .FEN(FEN[991]), .op(N2481_t1) );
fim FAN_N2484_0 ( .fault(fault), .net(N2484), .FEN(FEN[992]), .op(N2484_t0) );
fim FAN_N2484_1 ( .fault(fault), .net(N2484), .FEN(FEN[993]), .op(N2484_t1) );
fim FAN_N2417_0 ( .fault(fault), .net(N2417), .FEN(FEN[994]), .op(N2417_t0) );
fim FAN_N2417_1 ( .fault(fault), .net(N2417), .FEN(FEN[995]), .op(N2417_t1) );
fim FAN_N2417_2 ( .fault(fault), .net(N2417), .FEN(FEN[996]), .op(N2417_t2) );
fim FAN_N2421_0 ( .fault(fault), .net(N2421), .FEN(FEN[997]), .op(N2421_t0) );
fim FAN_N2421_1 ( .fault(fault), .net(N2421), .FEN(FEN[998]), .op(N2421_t1) );
fim FAN_N2421_2 ( .fault(fault), .net(N2421), .FEN(FEN[999]), .op(N2421_t2) );
fim FAN_N2425_0 ( .fault(fault), .net(N2425), .FEN(FEN[1000]), .op(N2425_t0) );
fim FAN_N2425_1 ( .fault(fault), .net(N2425), .FEN(FEN[1001]), .op(N2425_t1) );
fim FAN_N2493_0 ( .fault(fault), .net(N2493), .FEN(FEN[1002]), .op(N2493_t0) );
fim FAN_N2493_1 ( .fault(fault), .net(N2493), .FEN(FEN[1003]), .op(N2493_t1) );
fim FAN_N2440_0 ( .fault(fault), .net(N2440), .FEN(FEN[1004]), .op(N2440_t0) );
fim FAN_N2440_1 ( .fault(fault), .net(N2440), .FEN(FEN[1005]), .op(N2440_t1) );
fim FAN_N2443_0 ( .fault(fault), .net(N2443), .FEN(FEN[1006]), .op(N2443_t0) );
fim FAN_N2443_1 ( .fault(fault), .net(N2443), .FEN(FEN[1007]), .op(N2443_t1) );
fim FAN_N2446_0 ( .fault(fault), .net(N2446), .FEN(FEN[1008]), .op(N2446_t0) );
fim FAN_N2446_1 ( .fault(fault), .net(N2446), .FEN(FEN[1009]), .op(N2446_t1) );
fim FAN_N2449_0 ( .fault(fault), .net(N2449), .FEN(FEN[1010]), .op(N2449_t0) );
fim FAN_N2449_1 ( .fault(fault), .net(N2449), .FEN(FEN[1011]), .op(N2449_t1) );
fim FAN_N2457_0 ( .fault(fault), .net(N2457), .FEN(FEN[1012]), .op(N2457_t0) );
fim FAN_N2457_1 ( .fault(fault), .net(N2457), .FEN(FEN[1013]), .op(N2457_t1) );
fim FAN_N2460_0 ( .fault(fault), .net(N2460), .FEN(FEN[1014]), .op(N2460_t0) );
fim FAN_N2460_1 ( .fault(fault), .net(N2460), .FEN(FEN[1015]), .op(N2460_t1) );
fim FAN_N2463_0 ( .fault(fault), .net(N2463), .FEN(FEN[1016]), .op(N2463_t0) );
fim FAN_N2463_1 ( .fault(fault), .net(N2463), .FEN(FEN[1017]), .op(N2463_t1) );
fim FAN_N2466_0 ( .fault(fault), .net(N2466), .FEN(FEN[1018]), .op(N2466_t0) );
fim FAN_N2466_1 ( .fault(fault), .net(N2466), .FEN(FEN[1019]), .op(N2466_t1) );
fim FAN_N2469_0 ( .fault(fault), .net(N2469), .FEN(FEN[1020]), .op(N2469_t0) );
fim FAN_N2469_1 ( .fault(fault), .net(N2469), .FEN(FEN[1021]), .op(N2469_t1) );
fim FAN_N2487_0 ( .fault(fault), .net(N2487), .FEN(FEN[1022]), .op(N2487_t0) );
fim FAN_N2487_1 ( .fault(fault), .net(N2487), .FEN(FEN[1023]), .op(N2487_t1) );
fim FAN_N2490_0 ( .fault(fault), .net(N2490), .FEN(FEN[1024]), .op(N2490_t0) );
fim FAN_N2490_1 ( .fault(fault), .net(N2490), .FEN(FEN[1025]), .op(N2490_t1) );
fim FAN_N2534_0 ( .fault(fault), .net(N2534), .FEN(FEN[1026]), .op(N2534_t0) );
fim FAN_N2534_1 ( .fault(fault), .net(N2534), .FEN(FEN[1027]), .op(N2534_t1) );
fim FAN_N2531_0 ( .fault(fault), .net(N2531), .FEN(FEN[1028]), .op(N2531_t0) );
fim FAN_N2531_1 ( .fault(fault), .net(N2531), .FEN(FEN[1029]), .op(N2531_t1) );
fim FAN_N2537_0 ( .fault(fault), .net(N2537), .FEN(FEN[1030]), .op(N2537_t0) );
fim FAN_N2537_1 ( .fault(fault), .net(N2537), .FEN(FEN[1031]), .op(N2537_t1) );
fim FAN_N2540_0 ( .fault(fault), .net(N2540), .FEN(FEN[1032]), .op(N2540_t0) );
fim FAN_N2540_1 ( .fault(fault), .net(N2540), .FEN(FEN[1033]), .op(N2540_t1) );
fim FAN_N2638_0 ( .fault(fault), .net(N2638), .FEN(FEN[1034]), .op(N2638_t0) );
fim FAN_N2638_1 ( .fault(fault), .net(N2638), .FEN(FEN[1035]), .op(N2638_t1) );
fim FAN_N2638_2 ( .fault(fault), .net(N2638), .FEN(FEN[1036]), .op(N2638_t2) );
fim FAN_N2638_3 ( .fault(fault), .net(N2638), .FEN(FEN[1037]), .op(N2638_t3) );
fim FAN_N2613_0 ( .fault(fault), .net(N2613), .FEN(FEN[1038]), .op(N2613_t0) );
fim FAN_N2613_1 ( .fault(fault), .net(N2613), .FEN(FEN[1039]), .op(N2613_t1) );
fim FAN_N2613_2 ( .fault(fault), .net(N2613), .FEN(FEN[1040]), .op(N2613_t2) );
fim FAN_N2624_0 ( .fault(fault), .net(N2624), .FEN(FEN[1041]), .op(N2624_t0) );
fim FAN_N2624_1 ( .fault(fault), .net(N2624), .FEN(FEN[1042]), .op(N2624_t1) );
fim FAN_N2624_2 ( .fault(fault), .net(N2624), .FEN(FEN[1043]), .op(N2624_t2) );
fim FAN_N2646_0 ( .fault(fault), .net(N2646), .FEN(FEN[1044]), .op(N2646_t0) );
fim FAN_N2646_1 ( .fault(fault), .net(N2646), .FEN(FEN[1045]), .op(N2646_t1) );
fim FAN_N2646_2 ( .fault(fault), .net(N2646), .FEN(FEN[1046]), .op(N2646_t2) );
fim FAN_N2646_3 ( .fault(fault), .net(N2646), .FEN(FEN[1047]), .op(N2646_t3) );
fim FAN_N2603_0 ( .fault(fault), .net(N2603), .FEN(FEN[1048]), .op(N2603_t0) );
fim FAN_N2603_1 ( .fault(fault), .net(N2603), .FEN(FEN[1049]), .op(N2603_t1) );
fim FAN_N2603_2 ( .fault(fault), .net(N2603), .FEN(FEN[1050]), .op(N2603_t2) );
fim FAN_N2659_0 ( .fault(fault), .net(N2659), .FEN(FEN[1051]), .op(N2659_t0) );
fim FAN_N2659_1 ( .fault(fault), .net(N2659), .FEN(FEN[1052]), .op(N2659_t1) );
fim FAN_N2659_2 ( .fault(fault), .net(N2659), .FEN(FEN[1053]), .op(N2659_t2) );
fim FAN_N2687_0 ( .fault(fault), .net(N2687), .FEN(FEN[1054]), .op(N2687_t0) );
fim FAN_N2687_1 ( .fault(fault), .net(N2687), .FEN(FEN[1055]), .op(N2687_t1) );
fim FAN_N2690_0 ( .fault(fault), .net(N2690), .FEN(FEN[1056]), .op(N2690_t0) );
fim FAN_N2690_1 ( .fault(fault), .net(N2690), .FEN(FEN[1057]), .op(N2690_t1) );
fim FAN_N2684_0 ( .fault(fault), .net(N2684), .FEN(FEN[1058]), .op(N2684_t0) );
fim FAN_N2684_1 ( .fault(fault), .net(N2684), .FEN(FEN[1059]), .op(N2684_t1) );
fim FAN_N2681_0 ( .fault(fault), .net(N2681), .FEN(FEN[1060]), .op(N2681_t0) );
fim FAN_N2681_1 ( .fault(fault), .net(N2681), .FEN(FEN[1061]), .op(N2681_t1) );
fim FAN_N2703_0 ( .fault(fault), .net(N2703), .FEN(FEN[1062]), .op(N2703_t0) );
fim FAN_N2703_1 ( .fault(fault), .net(N2703), .FEN(FEN[1063]), .op(N2703_t1) );
fim FAN_N2729_0 ( .fault(fault), .net(N2729), .FEN(FEN[1064]), .op(N2729_t0) );
fim FAN_N2729_1 ( .fault(fault), .net(N2729), .FEN(FEN[1065]), .op(N2729_t1) );
fim FAN_N2729_2 ( .fault(fault), .net(N2729), .FEN(FEN[1066]), .op(N2729_t2) );
fim FAN_N2729_3 ( .fault(fault), .net(N2729), .FEN(FEN[1067]), .op(N2729_t3) );
fim FAN_N1037_0 ( .fault(fault), .net(N1037), .FEN(FEN[1068]), .op(N1037_t0) );
fim FAN_N1037_1 ( .fault(fault), .net(N1037), .FEN(FEN[1069]), .op(N1037_t1) );
fim FAN_N1037_2 ( .fault(fault), .net(N1037), .FEN(FEN[1070]), .op(N1037_t2) );
fim FAN_N1037_3 ( .fault(fault), .net(N1037), .FEN(FEN[1071]), .op(N1037_t3) );
fim FAN_N1070_0 ( .fault(fault), .net(N1070), .FEN(FEN[1072]), .op(N1070_t0) );
fim FAN_N1070_1 ( .fault(fault), .net(N1070), .FEN(FEN[1073]), .op(N1070_t1) );
fim FAN_N1070_2 ( .fault(fault), .net(N1070), .FEN(FEN[1074]), .op(N1070_t2) );
fim FAN_N1070_3 ( .fault(fault), .net(N1070), .FEN(FEN[1075]), .op(N1070_t3) );
fim FAN_N2738_0 ( .fault(fault), .net(N2738), .FEN(FEN[1076]), .op(N2738_t0) );
fim FAN_N2738_1 ( .fault(fault), .net(N2738), .FEN(FEN[1077]), .op(N2738_t1) );
fim FAN_N2738_2 ( .fault(fault), .net(N2738), .FEN(FEN[1078]), .op(N2738_t2) );
fim FAN_N2738_3 ( .fault(fault), .net(N2738), .FEN(FEN[1079]), .op(N2738_t3) );
fim FAN_N2817_0 ( .fault(fault), .net(N2817), .FEN(FEN[1080]), .op(N2817_t0) );
fim FAN_N2817_1 ( .fault(fault), .net(N2817), .FEN(FEN[1081]), .op(N2817_t1) );
fim FAN_N2841_0 ( .fault(fault), .net(N2841), .FEN(FEN[1082]), .op(N2841_t0) );
fim FAN_N2841_1 ( .fault(fault), .net(N2841), .FEN(FEN[1083]), .op(N2841_t1) );
fim FAN_N2826_0 ( .fault(fault), .net(N2826), .FEN(FEN[1084]), .op(N2826_t0) );
fim FAN_N2826_1 ( .fault(fault), .net(N2826), .FEN(FEN[1085]), .op(N2826_t1) );
fim FAN_N2796_0 ( .fault(fault), .net(N2796), .FEN(FEN[1086]), .op(N2796_t0) );
fim FAN_N2796_1 ( .fault(fault), .net(N2796), .FEN(FEN[1087]), .op(N2796_t1) );
fim FAN_N2796_2 ( .fault(fault), .net(N2796), .FEN(FEN[1088]), .op(N2796_t2) );
fim FAN_N2800_0 ( .fault(fault), .net(N2800), .FEN(FEN[1089]), .op(N2800_t0) );
fim FAN_N2800_1 ( .fault(fault), .net(N2800), .FEN(FEN[1090]), .op(N2800_t1) );
fim FAN_N2806_0 ( .fault(fault), .net(N2806), .FEN(FEN[1091]), .op(N2806_t0) );
fim FAN_N2806_1 ( .fault(fault), .net(N2806), .FEN(FEN[1092]), .op(N2806_t1) );
fim FAN_N2820_0 ( .fault(fault), .net(N2820), .FEN(FEN[1093]), .op(N2820_t0) );
fim FAN_N2820_1 ( .fault(fault), .net(N2820), .FEN(FEN[1094]), .op(N2820_t1) );
fim FAN_N2820_2 ( .fault(fault), .net(N2820), .FEN(FEN[1095]), .op(N2820_t2) );
fim FAN_N2820_3 ( .fault(fault), .net(N2820), .FEN(FEN[1096]), .op(N2820_t3) );
fim FAN_N2820_4 ( .fault(fault), .net(N2820), .FEN(FEN[1097]), .op(N2820_t4) );
fim FAN_N2831_0 ( .fault(fault), .net(N2831), .FEN(FEN[1098]), .op(N2831_t0) );
fim FAN_N2831_1 ( .fault(fault), .net(N2831), .FEN(FEN[1099]), .op(N2831_t1) );
fim FAN_N2831_2 ( .fault(fault), .net(N2831), .FEN(FEN[1100]), .op(N2831_t2) );
fim FAN_N2831_3 ( .fault(fault), .net(N2831), .FEN(FEN[1101]), .op(N2831_t3) );
fim FAN_N2831_4 ( .fault(fault), .net(N2831), .FEN(FEN[1102]), .op(N2831_t4) );
fim FAN_N2931_0 ( .fault(fault), .net(N2931), .FEN(FEN[1103]), .op(N2931_t0) );
fim FAN_N2931_1 ( .fault(fault), .net(N2931), .FEN(FEN[1104]), .op(N2931_t1) );
fim FAN_N2888_0 ( .fault(fault), .net(N2888), .FEN(FEN[1105]), .op(N2888_t0) );
fim FAN_N2888_1 ( .fault(fault), .net(N2888), .FEN(FEN[1106]), .op(N2888_t1) );
fim FAN_N2844_0 ( .fault(fault), .net(N2844), .FEN(FEN[1107]), .op(N2844_t0) );
fim FAN_N2844_1 ( .fault(fault), .net(N2844), .FEN(FEN[1108]), .op(N2844_t1) );
fim FAN_N2844_2 ( .fault(fault), .net(N2844), .FEN(FEN[1109]), .op(N2844_t2) );
fim FAN_N2844_3 ( .fault(fault), .net(N2844), .FEN(FEN[1110]), .op(N2844_t3) );
fim FAN_N2844_4 ( .fault(fault), .net(N2844), .FEN(FEN[1111]), .op(N2844_t4) );
fim FAN_N2854_0 ( .fault(fault), .net(N2854), .FEN(FEN[1112]), .op(N2854_t0) );
fim FAN_N2854_1 ( .fault(fault), .net(N2854), .FEN(FEN[1113]), .op(N2854_t1) );
fim FAN_N2854_2 ( .fault(fault), .net(N2854), .FEN(FEN[1114]), .op(N2854_t2) );
fim FAN_N2854_3 ( .fault(fault), .net(N2854), .FEN(FEN[1115]), .op(N2854_t3) );
fim FAN_N2859_0 ( .fault(fault), .net(N2859), .FEN(FEN[1116]), .op(N2859_t0) );
fim FAN_N2859_1 ( .fault(fault), .net(N2859), .FEN(FEN[1117]), .op(N2859_t1) );
fim FAN_N2859_2 ( .fault(fault), .net(N2859), .FEN(FEN[1118]), .op(N2859_t2) );
fim FAN_N2859_3 ( .fault(fault), .net(N2859), .FEN(FEN[1119]), .op(N2859_t3) );
fim FAN_N2859_4 ( .fault(fault), .net(N2859), .FEN(FEN[1120]), .op(N2859_t4) );
fim FAN_N2869_0 ( .fault(fault), .net(N2869), .FEN(FEN[1121]), .op(N2869_t0) );
fim FAN_N2869_1 ( .fault(fault), .net(N2869), .FEN(FEN[1122]), .op(N2869_t1) );
fim FAN_N2869_2 ( .fault(fault), .net(N2869), .FEN(FEN[1123]), .op(N2869_t2) );
fim FAN_N2869_3 ( .fault(fault), .net(N2869), .FEN(FEN[1124]), .op(N2869_t3) );
fim FAN_N2874_0 ( .fault(fault), .net(N2874), .FEN(FEN[1125]), .op(N2874_t0) );
fim FAN_N2874_1 ( .fault(fault), .net(N2874), .FEN(FEN[1126]), .op(N2874_t1) );
fim FAN_N2877_0 ( .fault(fault), .net(N2877), .FEN(FEN[1127]), .op(N2877_t0) );
fim FAN_N2877_1 ( .fault(fault), .net(N2877), .FEN(FEN[1128]), .op(N2877_t1) );
fim FAN_N2882_0 ( .fault(fault), .net(N2882), .FEN(FEN[1129]), .op(N2882_t0) );
fim FAN_N2882_1 ( .fault(fault), .net(N2882), .FEN(FEN[1130]), .op(N2882_t1) );
fim FAN_N2885_0 ( .fault(fault), .net(N2885), .FEN(FEN[1131]), .op(N2885_t0) );
fim FAN_N2885_1 ( .fault(fault), .net(N2885), .FEN(FEN[1132]), .op(N2885_t1) );
fim FAN_N1190_0 ( .fault(fault), .net(N1190), .FEN(FEN[1133]), .op(N1190_t0) );
fim FAN_N1190_1 ( .fault(fault), .net(N1190), .FEN(FEN[1134]), .op(N1190_t1) );
fim FAN_N1190_2 ( .fault(fault), .net(N1190), .FEN(FEN[1135]), .op(N1190_t2) );
fim FAN_N1190_3 ( .fault(fault), .net(N1190), .FEN(FEN[1136]), .op(N1190_t3) );
fim FAN_N2761_0 ( .fault(fault), .net(N2761), .FEN(FEN[1137]), .op(N2761_t0) );
fim FAN_N2761_1 ( .fault(fault), .net(N2761), .FEN(FEN[1138]), .op(N2761_t1) );
fim FAN_N2761_2 ( .fault(fault), .net(N2761), .FEN(FEN[1139]), .op(N2761_t2) );
fim FAN_N2761_3 ( .fault(fault), .net(N2761), .FEN(FEN[1140]), .op(N2761_t3) );
fim FAN_N1195_0 ( .fault(fault), .net(N1195), .FEN(FEN[1141]), .op(N1195_t0) );
fim FAN_N1195_1 ( .fault(fault), .net(N1195), .FEN(FEN[1142]), .op(N1195_t1) );
fim FAN_N1195_2 ( .fault(fault), .net(N1195), .FEN(FEN[1143]), .op(N1195_t2) );
fim FAN_N1195_3 ( .fault(fault), .net(N1195), .FEN(FEN[1144]), .op(N1195_t3) );
fim FAN_N2766_0 ( .fault(fault), .net(N2766), .FEN(FEN[1145]), .op(N2766_t0) );
fim FAN_N2766_1 ( .fault(fault), .net(N2766), .FEN(FEN[1146]), .op(N2766_t1) );
fim FAN_N2766_2 ( .fault(fault), .net(N2766), .FEN(FEN[1147]), .op(N2766_t2) );
fim FAN_N2766_3 ( .fault(fault), .net(N2766), .FEN(FEN[1148]), .op(N2766_t3) );
fim FAN_N2995_0 ( .fault(fault), .net(N2995), .FEN(FEN[1149]), .op(N2995_t0) );
fim FAN_N2995_1 ( .fault(fault), .net(N2995), .FEN(FEN[1150]), .op(N2995_t1) );
fim FAN_N2998_0 ( .fault(fault), .net(N2998), .FEN(FEN[1151]), .op(N2998_t0) );
fim FAN_N2998_1 ( .fault(fault), .net(N2998), .FEN(FEN[1152]), .op(N2998_t1) );
fim FAN_N3001_0 ( .fault(fault), .net(N3001), .FEN(FEN[1153]), .op(N3001_t0) );
fim FAN_N3001_1 ( .fault(fault), .net(N3001), .FEN(FEN[1154]), .op(N3001_t1) );
fim FAN_N3004_0 ( .fault(fault), .net(N3004), .FEN(FEN[1155]), .op(N3004_t0) );
fim FAN_N3004_1 ( .fault(fault), .net(N3004), .FEN(FEN[1156]), .op(N3004_t1) );
fim FAN_N2992_0 ( .fault(fault), .net(N2992), .FEN(FEN[1157]), .op(N2992_t0) );
fim FAN_N2992_1 ( .fault(fault), .net(N2992), .FEN(FEN[1158]), .op(N2992_t1) );
fim FAN_N2793_0 ( .fault(fault), .net(N2793), .FEN(FEN[1159]), .op(N2793_t0) );
fim FAN_N2793_1 ( .fault(fault), .net(N2793), .FEN(FEN[1160]), .op(N2793_t1) );
fim FAN_N2803_0 ( .fault(fault), .net(N2803), .FEN(FEN[1161]), .op(N2803_t0) );
fim FAN_N2803_1 ( .fault(fault), .net(N2803), .FEN(FEN[1162]), .op(N2803_t1) );
fim FAN_N2621_0 ( .fault(fault), .net(N2621), .FEN(FEN[1163]), .op(N2621_t0) );
fim FAN_N2621_1 ( .fault(fault), .net(N2621), .FEN(FEN[1164]), .op(N2621_t1) );
fim FAN_N3076_0 ( .fault(fault), .net(N3076), .FEN(FEN[1165]), .op(N3076_t0) );
fim FAN_N3076_1 ( .fault(fault), .net(N3076), .FEN(FEN[1166]), .op(N3076_t1) );
fim FAN_N3030_0 ( .fault(fault), .net(N3030), .FEN(FEN[1167]), .op(N3030_t0) );
fim FAN_N3030_1 ( .fault(fault), .net(N3030), .FEN(FEN[1168]), .op(N3030_t1) );
fim FAN_N3030_2 ( .fault(fault), .net(N3030), .FEN(FEN[1169]), .op(N3030_t2) );
fim FAN_N3030_3 ( .fault(fault), .net(N3030), .FEN(FEN[1170]), .op(N3030_t3) );
fim FAN_N3039_0 ( .fault(fault), .net(N3039), .FEN(FEN[1171]), .op(N3039_t0) );
fim FAN_N3039_1 ( .fault(fault), .net(N3039), .FEN(FEN[1172]), .op(N3039_t1) );
fim FAN_N3039_2 ( .fault(fault), .net(N3039), .FEN(FEN[1173]), .op(N3039_t2) );
fim FAN_N3039_3 ( .fault(fault), .net(N3039), .FEN(FEN[1174]), .op(N3039_t3) );
fim FAN_N3050_0 ( .fault(fault), .net(N3050), .FEN(FEN[1175]), .op(N3050_t0) );
fim FAN_N3050_1 ( .fault(fault), .net(N3050), .FEN(FEN[1176]), .op(N3050_t1) );
fim FAN_N3061_0 ( .fault(fault), .net(N3061), .FEN(FEN[1177]), .op(N3061_t0) );
fim FAN_N3061_1 ( .fault(fault), .net(N3061), .FEN(FEN[1178]), .op(N3061_t1) );
fim FAN_N2981_0 ( .fault(fault), .net(N2981), .FEN(FEN[1179]), .op(N2981_t0) );
fim FAN_N2981_1 ( .fault(fault), .net(N2981), .FEN(FEN[1180]), .op(N2981_t1) );
fim FAN_N2978_0 ( .fault(fault), .net(N2978), .FEN(FEN[1181]), .op(N2978_t0) );
fim FAN_N2978_1 ( .fault(fault), .net(N2978), .FEN(FEN[1182]), .op(N2978_t1) );
fim FAN_N2975_0 ( .fault(fault), .net(N2975), .FEN(FEN[1183]), .op(N2975_t0) );
fim FAN_N2975_1 ( .fault(fault), .net(N2975), .FEN(FEN[1184]), .op(N2975_t1) );
fim FAN_N2972_0 ( .fault(fault), .net(N2972), .FEN(FEN[1185]), .op(N2972_t0) );
fim FAN_N2972_1 ( .fault(fault), .net(N2972), .FEN(FEN[1186]), .op(N2972_t1) );
fim FAN_N2989_0 ( .fault(fault), .net(N2989), .FEN(FEN[1187]), .op(N2989_t0) );
fim FAN_N2989_1 ( .fault(fault), .net(N2989), .FEN(FEN[1188]), .op(N2989_t1) );
fim FAN_N2986_0 ( .fault(fault), .net(N2986), .FEN(FEN[1189]), .op(N2986_t0) );
fim FAN_N2986_1 ( .fault(fault), .net(N2986), .FEN(FEN[1190]), .op(N2986_t1) );
fim FAN_N3025_0 ( .fault(fault), .net(N3025), .FEN(FEN[1191]), .op(N3025_t0) );
fim FAN_N3025_1 ( .fault(fault), .net(N3025), .FEN(FEN[1192]), .op(N3025_t1) );
fim FAN_N3022_0 ( .fault(fault), .net(N3022), .FEN(FEN[1193]), .op(N3022_t0) );
fim FAN_N3022_1 ( .fault(fault), .net(N3022), .FEN(FEN[1194]), .op(N3022_t1) );
fim FAN_N3019_0 ( .fault(fault), .net(N3019), .FEN(FEN[1195]), .op(N3019_t0) );
fim FAN_N3019_1 ( .fault(fault), .net(N3019), .FEN(FEN[1196]), .op(N3019_t1) );
fim FAN_N3016_0 ( .fault(fault), .net(N3016), .FEN(FEN[1197]), .op(N3016_t0) );
fim FAN_N3016_1 ( .fault(fault), .net(N3016), .FEN(FEN[1198]), .op(N3016_t1) );
fim FAN_N3013_0 ( .fault(fault), .net(N3013), .FEN(FEN[1199]), .op(N3013_t0) );
fim FAN_N3013_1 ( .fault(fault), .net(N3013), .FEN(FEN[1200]), .op(N3013_t1) );
fim FAN_N3010_0 ( .fault(fault), .net(N3010), .FEN(FEN[1201]), .op(N3010_t0) );
fim FAN_N3010_1 ( .fault(fault), .net(N3010), .FEN(FEN[1202]), .op(N3010_t1) );
fim FAN_N3180_0 ( .fault(fault), .net(N3180), .FEN(FEN[1203]), .op(N3180_t0) );
fim FAN_N3180_1 ( .fault(fault), .net(N3180), .FEN(FEN[1204]), .op(N3180_t1) );
fim FAN_N3152_0 ( .fault(fault), .net(N3152), .FEN(FEN[1205]), .op(N3152_t0) );
fim FAN_N3152_1 ( .fault(fault), .net(N3152), .FEN(FEN[1206]), .op(N3152_t1) );
fim FAN_N3149_0 ( .fault(fault), .net(N3149), .FEN(FEN[1207]), .op(N3149_t0) );
fim FAN_N3149_1 ( .fault(fault), .net(N3149), .FEN(FEN[1208]), .op(N3149_t1) );
fim FAN_N3146_0 ( .fault(fault), .net(N3146), .FEN(FEN[1209]), .op(N3146_t0) );
fim FAN_N3146_1 ( .fault(fault), .net(N3146), .FEN(FEN[1210]), .op(N3146_t1) );
fim FAN_N3143_0 ( .fault(fault), .net(N3143), .FEN(FEN[1211]), .op(N3143_t0) );
fim FAN_N3143_1 ( .fault(fault), .net(N3143), .FEN(FEN[1212]), .op(N3143_t1) );
fim FAN_N3140_0 ( .fault(fault), .net(N3140), .FEN(FEN[1213]), .op(N3140_t0) );
fim FAN_N3140_1 ( .fault(fault), .net(N3140), .FEN(FEN[1214]), .op(N3140_t1) );
fim FAN_N3137_0 ( .fault(fault), .net(N3137), .FEN(FEN[1215]), .op(N3137_t0) );
fim FAN_N3137_1 ( .fault(fault), .net(N3137), .FEN(FEN[1216]), .op(N3137_t1) );
fim FAN_N3172_0 ( .fault(fault), .net(N3172), .FEN(FEN[1217]), .op(N3172_t0) );
fim FAN_N3172_1 ( .fault(fault), .net(N3172), .FEN(FEN[1218]), .op(N3172_t1) );
fim FAN_N3169_0 ( .fault(fault), .net(N3169), .FEN(FEN[1219]), .op(N3169_t0) );
fim FAN_N3169_1 ( .fault(fault), .net(N3169), .FEN(FEN[1220]), .op(N3169_t1) );
fim FAN_N3166_0 ( .fault(fault), .net(N3166), .FEN(FEN[1221]), .op(N3166_t0) );
fim FAN_N3166_1 ( .fault(fault), .net(N3166), .FEN(FEN[1222]), .op(N3166_t1) );
fim FAN_N3163_0 ( .fault(fault), .net(N3163), .FEN(FEN[1223]), .op(N3163_t0) );
fim FAN_N3163_1 ( .fault(fault), .net(N3163), .FEN(FEN[1224]), .op(N3163_t1) );
fim FAN_N3160_0 ( .fault(fault), .net(N3160), .FEN(FEN[1225]), .op(N3160_t0) );
fim FAN_N3160_1 ( .fault(fault), .net(N3160), .FEN(FEN[1226]), .op(N3160_t1) );
fim FAN_N3157_0 ( .fault(fault), .net(N3157), .FEN(FEN[1227]), .op(N3157_t0) );
fim FAN_N3157_1 ( .fault(fault), .net(N3157), .FEN(FEN[1228]), .op(N3157_t1) );
fim FAN_N3091_0 ( .fault(fault), .net(N3091), .FEN(FEN[1229]), .op(N3091_t0) );
fim FAN_N3091_1 ( .fault(fault), .net(N3091), .FEN(FEN[1230]), .op(N3091_t1) );
fim FAN_N3088_0 ( .fault(fault), .net(N3088), .FEN(FEN[1231]), .op(N3088_t0) );
fim FAN_N3088_1 ( .fault(fault), .net(N3088), .FEN(FEN[1232]), .op(N3088_t1) );
fim FAN_N3113_0 ( .fault(fault), .net(N3113), .FEN(FEN[1233]), .op(N3113_t0) );
fim FAN_N3113_1 ( .fault(fault), .net(N3113), .FEN(FEN[1234]), .op(N3113_t1) );
fim FAN_N3110_0 ( .fault(fault), .net(N3110), .FEN(FEN[1235]), .op(N3110_t0) );
fim FAN_N3110_1 ( .fault(fault), .net(N3110), .FEN(FEN[1236]), .op(N3110_t1) );
fim FAN_N3238_0 ( .fault(fault), .net(N3238), .FEN(FEN[1237]), .op(N3238_t0) );
fim FAN_N3238_1 ( .fault(fault), .net(N3238), .FEN(FEN[1238]), .op(N3238_t1) );
fim FAN_N3241_0 ( .fault(fault), .net(N3241), .FEN(FEN[1239]), .op(N3241_t0) );
fim FAN_N3241_1 ( .fault(fault), .net(N3241), .FEN(FEN[1240]), .op(N3241_t1) );
fim FAN_N3244_0 ( .fault(fault), .net(N3244), .FEN(FEN[1241]), .op(N3244_t0) );
fim FAN_N3244_1 ( .fault(fault), .net(N3244), .FEN(FEN[1242]), .op(N3244_t1) );
fim FAN_N3247_0 ( .fault(fault), .net(N3247), .FEN(FEN[1243]), .op(N3247_t0) );
fim FAN_N3247_1 ( .fault(fault), .net(N3247), .FEN(FEN[1244]), .op(N3247_t1) );
fim FAN_N3250_0 ( .fault(fault), .net(N3250), .FEN(FEN[1245]), .op(N3250_t0) );
fim FAN_N3250_1 ( .fault(fault), .net(N3250), .FEN(FEN[1246]), .op(N3250_t1) );
fim FAN_N3253_0 ( .fault(fault), .net(N3253), .FEN(FEN[1247]), .op(N3253_t0) );
fim FAN_N3253_1 ( .fault(fault), .net(N3253), .FEN(FEN[1248]), .op(N3253_t1) );
fim FAN_N3256_0 ( .fault(fault), .net(N3256), .FEN(FEN[1249]), .op(N3256_t0) );
fim FAN_N3256_1 ( .fault(fault), .net(N3256), .FEN(FEN[1250]), .op(N3256_t1) );
fim FAN_N3259_0 ( .fault(fault), .net(N3259), .FEN(FEN[1251]), .op(N3259_t0) );
fim FAN_N3259_1 ( .fault(fault), .net(N3259), .FEN(FEN[1252]), .op(N3259_t1) );
fim FAN_N3262_0 ( .fault(fault), .net(N3262), .FEN(FEN[1253]), .op(N3262_t0) );
fim FAN_N3262_1 ( .fault(fault), .net(N3262), .FEN(FEN[1254]), .op(N3262_t1) );
fim FAN_N3265_0 ( .fault(fault), .net(N3265), .FEN(FEN[1255]), .op(N3265_t0) );
fim FAN_N3265_1 ( .fault(fault), .net(N3265), .FEN(FEN[1256]), .op(N3265_t1) );
fim FAN_N3268_0 ( .fault(fault), .net(N3268), .FEN(FEN[1257]), .op(N3268_t0) );
fim FAN_N3268_1 ( .fault(fault), .net(N3268), .FEN(FEN[1258]), .op(N3268_t1) );
fim FAN_N3271_0 ( .fault(fault), .net(N3271), .FEN(FEN[1259]), .op(N3271_t0) );
fim FAN_N3271_1 ( .fault(fault), .net(N3271), .FEN(FEN[1260]), .op(N3271_t1) );
fim FAN_N3274_0 ( .fault(fault), .net(N3274), .FEN(FEN[1261]), .op(N3274_t0) );
fim FAN_N3274_1 ( .fault(fault), .net(N3274), .FEN(FEN[1262]), .op(N3274_t1) );
fim FAN_N3277_0 ( .fault(fault), .net(N3277), .FEN(FEN[1263]), .op(N3277_t0) );
fim FAN_N3277_1 ( .fault(fault), .net(N3277), .FEN(FEN[1264]), .op(N3277_t1) );
fim FAN_N3318_0 ( .fault(fault), .net(N3318), .FEN(FEN[1265]), .op(N3318_t0) );
fim FAN_N3318_1 ( .fault(fault), .net(N3318), .FEN(FEN[1266]), .op(N3318_t1) );
fim FAN_N3315_0 ( .fault(fault), .net(N3315), .FEN(FEN[1267]), .op(N3315_t0) );
fim FAN_N3315_1 ( .fault(fault), .net(N3315), .FEN(FEN[1268]), .op(N3315_t1) );
fim FAN_N3340_0 ( .fault(fault), .net(N3340), .FEN(FEN[1269]), .op(N3340_t0) );
fim FAN_N3340_1 ( .fault(fault), .net(N3340), .FEN(FEN[1270]), .op(N3340_t1) );
fim FAN_N3344_0 ( .fault(fault), .net(N3344), .FEN(FEN[1271]), .op(N3344_t0) );
fim FAN_N3344_1 ( .fault(fault), .net(N3344), .FEN(FEN[1272]), .op(N3344_t1) );
fim FAN_N3348_0 ( .fault(fault), .net(N3348), .FEN(FEN[1273]), .op(N3348_t0) );
fim FAN_N3348_1 ( .fault(fault), .net(N3348), .FEN(FEN[1274]), .op(N3348_t1) );
fim FAN_N3352_0 ( .fault(fault), .net(N3352), .FEN(FEN[1275]), .op(N3352_t0) );
fim FAN_N3352_1 ( .fault(fault), .net(N3352), .FEN(FEN[1276]), .op(N3352_t1) );
fim FAN_N3356_0 ( .fault(fault), .net(N3356), .FEN(FEN[1277]), .op(N3356_t0) );
fim FAN_N3356_1 ( .fault(fault), .net(N3356), .FEN(FEN[1278]), .op(N3356_t1) );
fim FAN_N3360_0 ( .fault(fault), .net(N3360), .FEN(FEN[1279]), .op(N3360_t0) );
fim FAN_N3360_1 ( .fault(fault), .net(N3360), .FEN(FEN[1280]), .op(N3360_t1) );
fim FAN_N3364_0 ( .fault(fault), .net(N3364), .FEN(FEN[1281]), .op(N3364_t0) );
fim FAN_N3364_1 ( .fault(fault), .net(N3364), .FEN(FEN[1282]), .op(N3364_t1) );
fim FAN_N3367_0 ( .fault(fault), .net(N3367), .FEN(FEN[1283]), .op(N3367_t0) );
fim FAN_N3367_1 ( .fault(fault), .net(N3367), .FEN(FEN[1284]), .op(N3367_t1) );
fim FAN_N3321_0 ( .fault(fault), .net(N3321), .FEN(FEN[1285]), .op(N3321_t0) );
fim FAN_N3321_1 ( .fault(fault), .net(N3321), .FEN(FEN[1286]), .op(N3321_t1) );
fim FAN_N3327_0 ( .fault(fault), .net(N3327), .FEN(FEN[1287]), .op(N3327_t0) );
fim FAN_N3327_1 ( .fault(fault), .net(N3327), .FEN(FEN[1288]), .op(N3327_t1) );
fim FAN_N3324_0 ( .fault(fault), .net(N3324), .FEN(FEN[1289]), .op(N3324_t0) );
fim FAN_N3324_1 ( .fault(fault), .net(N3324), .FEN(FEN[1290]), .op(N3324_t1) );
fim FAN_N3370_0 ( .fault(fault), .net(N3370), .FEN(FEN[1291]), .op(N3370_t0) );
fim FAN_N3370_1 ( .fault(fault), .net(N3370), .FEN(FEN[1292]), .op(N3370_t1) );
fim FAN_N3374_0 ( .fault(fault), .net(N3374), .FEN(FEN[1293]), .op(N3374_t0) );
fim FAN_N3374_1 ( .fault(fault), .net(N3374), .FEN(FEN[1294]), .op(N3374_t1) );
fim FAN_N3378_0 ( .fault(fault), .net(N3378), .FEN(FEN[1295]), .op(N3378_t0) );
fim FAN_N3378_1 ( .fault(fault), .net(N3378), .FEN(FEN[1296]), .op(N3378_t1) );
fim FAN_N3382_0 ( .fault(fault), .net(N3382), .FEN(FEN[1297]), .op(N3382_t0) );
fim FAN_N3382_1 ( .fault(fault), .net(N3382), .FEN(FEN[1298]), .op(N3382_t1) );
fim FAN_N3386_0 ( .fault(fault), .net(N3386), .FEN(FEN[1299]), .op(N3386_t0) );
fim FAN_N3386_1 ( .fault(fault), .net(N3386), .FEN(FEN[1300]), .op(N3386_t1) );
fim FAN_N3390_0 ( .fault(fault), .net(N3390), .FEN(FEN[1301]), .op(N3390_t0) );
fim FAN_N3390_1 ( .fault(fault), .net(N3390), .FEN(FEN[1302]), .op(N3390_t1) );
fim FAN_N3394_0 ( .fault(fault), .net(N3394), .FEN(FEN[1303]), .op(N3394_t0) );
fim FAN_N3394_1 ( .fault(fault), .net(N3394), .FEN(FEN[1304]), .op(N3394_t1) );
fim FAN_N3397_0 ( .fault(fault), .net(N3397), .FEN(FEN[1305]), .op(N3397_t0) );
fim FAN_N3397_1 ( .fault(fault), .net(N3397), .FEN(FEN[1306]), .op(N3397_t1) );
fim FAN_N3330_0 ( .fault(fault), .net(N3330), .FEN(FEN[1307]), .op(N3330_t0) );
fim FAN_N3330_1 ( .fault(fault), .net(N3330), .FEN(FEN[1308]), .op(N3330_t1) );
fim FAN_N3453_0 ( .fault(fault), .net(N3453), .FEN(FEN[1309]), .op(N3453_t0) );
fim FAN_N3453_1 ( .fault(fault), .net(N3453), .FEN(FEN[1310]), .op(N3453_t1) );
fim FAN_N3450_0 ( .fault(fault), .net(N3450), .FEN(FEN[1311]), .op(N3450_t0) );
fim FAN_N3450_1 ( .fault(fault), .net(N3450), .FEN(FEN[1312]), .op(N3450_t1) );
fim FAN_N3459_0 ( .fault(fault), .net(N3459), .FEN(FEN[1313]), .op(N3459_t0) );
fim FAN_N3459_1 ( .fault(fault), .net(N3459), .FEN(FEN[1314]), .op(N3459_t1) );
fim FAN_N3456_0 ( .fault(fault), .net(N3456), .FEN(FEN[1315]), .op(N3456_t0) );
fim FAN_N3456_1 ( .fault(fault), .net(N3456), .FEN(FEN[1316]), .op(N3456_t1) );
fim FAN_N3522_0 ( .fault(fault), .net(N3522), .FEN(FEN[1317]), .op(N3522_t0) );
fim FAN_N3522_1 ( .fault(fault), .net(N3522), .FEN(FEN[1318]), .op(N3522_t1) );
fim FAN_N3525_0 ( .fault(fault), .net(N3525), .FEN(FEN[1319]), .op(N3525_t0) );
fim FAN_N3525_1 ( .fault(fault), .net(N3525), .FEN(FEN[1320]), .op(N3525_t1) );
fim FAN_N3528_0 ( .fault(fault), .net(N3528), .FEN(FEN[1321]), .op(N3528_t0) );
fim FAN_N3528_1 ( .fault(fault), .net(N3528), .FEN(FEN[1322]), .op(N3528_t1) );
fim FAN_N3531_0 ( .fault(fault), .net(N3531), .FEN(FEN[1323]), .op(N3531_t0) );
fim FAN_N3531_1 ( .fault(fault), .net(N3531), .FEN(FEN[1324]), .op(N3531_t1) );
fim FAN_N800_0 ( .fault(fault), .net(N800), .FEN(FEN[1325]), .op(N800_t0) );
fim FAN_N800_1 ( .fault(fault), .net(N800), .FEN(FEN[1326]), .op(N800_t1) );
fim FAN_N3534_0 ( .fault(fault), .net(N3534), .FEN(FEN[1327]), .op(N3534_t0) );
fim FAN_N3534_1 ( .fault(fault), .net(N3534), .FEN(FEN[1328]), .op(N3534_t1) );
fim FAN_N3537_0 ( .fault(fault), .net(N3537), .FEN(FEN[1329]), .op(N3537_t0) );
fim FAN_N3537_1 ( .fault(fault), .net(N3537), .FEN(FEN[1330]), .op(N3537_t1) );
fim FAN_N3540_0 ( .fault(fault), .net(N3540), .FEN(FEN[1331]), .op(N3540_t0) );
fim FAN_N3540_1 ( .fault(fault), .net(N3540), .FEN(FEN[1332]), .op(N3540_t1) );
fim FAN_N3543_0 ( .fault(fault), .net(N3543), .FEN(FEN[1333]), .op(N3543_t0) );
fim FAN_N3543_1 ( .fault(fault), .net(N3543), .FEN(FEN[1334]), .op(N3543_t1) );
fim FAN_N3600_0 ( .fault(fault), .net(N3600), .FEN(FEN[1335]), .op(N3600_t0) );
fim FAN_N3600_1 ( .fault(fault), .net(N3600), .FEN(FEN[1336]), .op(N3600_t1) );
fim FAN_N3576_0 ( .fault(fault), .net(N3576), .FEN(FEN[1337]), .op(N3576_t0) );
fim FAN_N3576_1 ( .fault(fault), .net(N3576), .FEN(FEN[1338]), .op(N3576_t1) );
fim FAN_N3579_0 ( .fault(fault), .net(N3579), .FEN(FEN[1339]), .op(N3579_t0) );
fim FAN_N3579_1 ( .fault(fault), .net(N3579), .FEN(FEN[1340]), .op(N3579_t1) );
fim FAN_N3585_0 ( .fault(fault), .net(N3585), .FEN(FEN[1341]), .op(N3585_t0) );
fim FAN_N3585_1 ( .fault(fault), .net(N3585), .FEN(FEN[1342]), .op(N3585_t1) );
fim FAN_N3588_0 ( .fault(fault), .net(N3588), .FEN(FEN[1343]), .op(N3588_t0) );
fim FAN_N3588_1 ( .fault(fault), .net(N3588), .FEN(FEN[1344]), .op(N3588_t1) );
fim FAN_N3608_0 ( .fault(fault), .net(N3608), .FEN(FEN[1345]), .op(N3608_t0) );
fim FAN_N3608_1 ( .fault(fault), .net(N3608), .FEN(FEN[1346]), .op(N3608_t1) );
fim FAN_N3608_2 ( .fault(fault), .net(N3608), .FEN(FEN[1347]), .op(N3608_t2) );
fim FAN_N3612_0 ( .fault(fault), .net(N3612), .FEN(FEN[1348]), .op(N3612_t0) );
fim FAN_N3612_1 ( .fault(fault), .net(N3612), .FEN(FEN[1349]), .op(N3612_t1) );
fim FAN_N3603_0 ( .fault(fault), .net(N3603), .FEN(FEN[1350]), .op(N3603_t0) );
fim FAN_N3603_1 ( .fault(fault), .net(N3603), .FEN(FEN[1351]), .op(N3603_t1) );
fim FAN_N3603_2 ( .fault(fault), .net(N3603), .FEN(FEN[1352]), .op(N3603_t2) );
fim FAN_N3603_3 ( .fault(fault), .net(N3603), .FEN(FEN[1353]), .op(N3603_t3) );
fim FAN_N3616_0 ( .fault(fault), .net(N3616), .FEN(FEN[1354]), .op(N3616_t0) );
fim FAN_N3616_1 ( .fault(fault), .net(N3616), .FEN(FEN[1355]), .op(N3616_t1) );
fim FAN_N3616_2 ( .fault(fault), .net(N3616), .FEN(FEN[1356]), .op(N3616_t2) );
fim FAN_N3616_3 ( .fault(fault), .net(N3616), .FEN(FEN[1357]), .op(N3616_t3) );
fim FAN_N3616_4 ( .fault(fault), .net(N3616), .FEN(FEN[1358]), .op(N3616_t4) );
fim FAN_N3622_0 ( .fault(fault), .net(N3622), .FEN(FEN[1359]), .op(N3622_t0) );
fim FAN_N3622_1 ( .fault(fault), .net(N3622), .FEN(FEN[1360]), .op(N3622_t1) );
fim FAN_N3622_2 ( .fault(fault), .net(N3622), .FEN(FEN[1361]), .op(N3622_t2) );
fim FAN_N3622_3 ( .fault(fault), .net(N3622), .FEN(FEN[1362]), .op(N3622_t3) );
fim FAN_N3640_0 ( .fault(fault), .net(N3640), .FEN(FEN[1363]), .op(N3640_t0) );
fim FAN_N3640_1 ( .fault(fault), .net(N3640), .FEN(FEN[1364]), .op(N3640_t1) );
fim FAN_N3640_2 ( .fault(fault), .net(N3640), .FEN(FEN[1365]), .op(N3640_t2) );
fim FAN_N3644_0 ( .fault(fault), .net(N3644), .FEN(FEN[1366]), .op(N3644_t0) );
fim FAN_N3644_1 ( .fault(fault), .net(N3644), .FEN(FEN[1367]), .op(N3644_t1) );
fim FAN_N3635_0 ( .fault(fault), .net(N3635), .FEN(FEN[1368]), .op(N3635_t0) );
fim FAN_N3635_1 ( .fault(fault), .net(N3635), .FEN(FEN[1369]), .op(N3635_t1) );
fim FAN_N3635_2 ( .fault(fault), .net(N3635), .FEN(FEN[1370]), .op(N3635_t2) );
fim FAN_N3635_3 ( .fault(fault), .net(N3635), .FEN(FEN[1371]), .op(N3635_t3) );
fim FAN_N3648_0 ( .fault(fault), .net(N3648), .FEN(FEN[1372]), .op(N3648_t0) );
fim FAN_N3648_1 ( .fault(fault), .net(N3648), .FEN(FEN[1373]), .op(N3648_t1) );
fim FAN_N3648_2 ( .fault(fault), .net(N3648), .FEN(FEN[1374]), .op(N3648_t2) );
fim FAN_N3648_3 ( .fault(fault), .net(N3648), .FEN(FEN[1375]), .op(N3648_t3) );
fim FAN_N3648_4 ( .fault(fault), .net(N3648), .FEN(FEN[1376]), .op(N3648_t4) );
fim FAN_N3654_0 ( .fault(fault), .net(N3654), .FEN(FEN[1377]), .op(N3654_t0) );
fim FAN_N3654_1 ( .fault(fault), .net(N3654), .FEN(FEN[1378]), .op(N3654_t1) );
fim FAN_N3654_2 ( .fault(fault), .net(N3654), .FEN(FEN[1379]), .op(N3654_t2) );
fim FAN_N3654_3 ( .fault(fault), .net(N3654), .FEN(FEN[1380]), .op(N3654_t3) );
fim FAN_N3723_0 ( .fault(fault), .net(N3723), .FEN(FEN[1381]), .op(N3723_t0) );
fim FAN_N3723_1 ( .fault(fault), .net(N3723), .FEN(FEN[1382]), .op(N3723_t1) );
fim FAN_N3737_0 ( .fault(fault), .net(N3737), .FEN(FEN[1383]), .op(N3737_t0) );
fim FAN_N3737_1 ( .fault(fault), .net(N3737), .FEN(FEN[1384]), .op(N3737_t1) );
fim FAN_N3780_0 ( .fault(fault), .net(N3780), .FEN(FEN[1385]), .op(N3780_t0) );
fim FAN_N3780_1 ( .fault(fault), .net(N3780), .FEN(FEN[1386]), .op(N3780_t1) );
fim FAN_N3762_0 ( .fault(fault), .net(N3762), .FEN(FEN[1387]), .op(N3762_t0) );
fim FAN_N3762_1 ( .fault(fault), .net(N3762), .FEN(FEN[1388]), .op(N3762_t1) );
fim FAN_N3754_0 ( .fault(fault), .net(N3754), .FEN(FEN[1389]), .op(N3754_t0) );
fim FAN_N3754_1 ( .fault(fault), .net(N3754), .FEN(FEN[1390]), .op(N3754_t1) );
fim FAN_N3754_2 ( .fault(fault), .net(N3754), .FEN(FEN[1391]), .op(N3754_t2) );
fim FAN_N3758_0 ( .fault(fault), .net(N3758), .FEN(FEN[1392]), .op(N3758_t0) );
fim FAN_N3758_1 ( .fault(fault), .net(N3758), .FEN(FEN[1393]), .op(N3758_t1) );
fim FAN_N3790_0 ( .fault(fault), .net(N3790), .FEN(FEN[1394]), .op(N3790_t0) );
fim FAN_N3790_1 ( .fault(fault), .net(N3790), .FEN(FEN[1395]), .op(N3790_t1) );
fim FAN_N3775_0 ( .fault(fault), .net(N3775), .FEN(FEN[1396]), .op(N3775_t0) );
fim FAN_N3775_1 ( .fault(fault), .net(N3775), .FEN(FEN[1397]), .op(N3775_t1) );
fim FAN_N3767_0 ( .fault(fault), .net(N3767), .FEN(FEN[1398]), .op(N3767_t0) );
fim FAN_N3767_1 ( .fault(fault), .net(N3767), .FEN(FEN[1399]), .op(N3767_t1) );
fim FAN_N3767_2 ( .fault(fault), .net(N3767), .FEN(FEN[1400]), .op(N3767_t2) );
fim FAN_N3771_0 ( .fault(fault), .net(N3771), .FEN(FEN[1401]), .op(N3771_t0) );
fim FAN_N3771_1 ( .fault(fault), .net(N3771), .FEN(FEN[1402]), .op(N3771_t1) );
fim FAN_N3823_0 ( .fault(fault), .net(N3823), .FEN(FEN[1403]), .op(N3823_t0) );
fim FAN_N3823_1 ( .fault(fault), .net(N3823), .FEN(FEN[1404]), .op(N3823_t1) );
fim FAN_N3827_0 ( .fault(fault), .net(N3827), .FEN(FEN[1405]), .op(N3827_t0) );
fim FAN_N3827_1 ( .fault(fault), .net(N3827), .FEN(FEN[1406]), .op(N3827_t1) );
fim FAN_N3843_0 ( .fault(fault), .net(N3843), .FEN(FEN[1407]), .op(N3843_t0) );
fim FAN_N3843_1 ( .fault(fault), .net(N3843), .FEN(FEN[1408]), .op(N3843_t1) );
fim FAN_N3843_2 ( .fault(fault), .net(N3843), .FEN(FEN[1409]), .op(N3843_t2) );
fim FAN_N3840_0 ( .fault(fault), .net(N3840), .FEN(FEN[1410]), .op(N3840_t0) );
fim FAN_N3840_1 ( .fault(fault), .net(N3840), .FEN(FEN[1411]), .op(N3840_t1) );
fim FAN_N3852_0 ( .fault(fault), .net(N3852), .FEN(FEN[1412]), .op(N3852_t0) );
fim FAN_N3852_1 ( .fault(fault), .net(N3852), .FEN(FEN[1413]), .op(N3852_t1) );
fim FAN_N3859_0 ( .fault(fault), .net(N3859), .FEN(FEN[1414]), .op(N3859_t0) );
fim FAN_N3859_1 ( .fault(fault), .net(N3859), .FEN(FEN[1415]), .op(N3859_t1) );
fim FAN_N3864_0 ( .fault(fault), .net(N3864), .FEN(FEN[1416]), .op(N3864_t0) );
fim FAN_N3864_1 ( .fault(fault), .net(N3864), .FEN(FEN[1417]), .op(N3864_t1) );
fim FAN_N3870_0 ( .fault(fault), .net(N3870), .FEN(FEN[1418]), .op(N3870_t0) );
fim FAN_N3870_1 ( .fault(fault), .net(N3870), .FEN(FEN[1419]), .op(N3870_t1) );
fim FAN_N3877_0 ( .fault(fault), .net(N3877), .FEN(FEN[1420]), .op(N3877_t0) );
fim FAN_N3877_1 ( .fault(fault), .net(N3877), .FEN(FEN[1421]), .op(N3877_t1) );
initial begin
    FEN <= {1421'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {1421'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,1421'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,1421'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN <= {FEN[1420:0], FEN[1421]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
// EndFaultModel

//Anchor
buf BUFF1_1 (N398, N219_t0);
buf BUFF1_2 (N400, N219_t1);
buf BUFF1_3 (N401, N219_t2);
and AND2_4 (N405, N1_t, N3_t);
not NOT1_5 (N408, N230_t);
buf BUFF1_6 (N419, N253_t0);
buf BUFF1_7 (N420, N253_t1);
not NOT1_8 (N425, N262_t);
buf BUFF1_9 (N456, N290_t0);
buf BUFF1_10 (N457, N290_t1);
buf BUFF1_11 (N458, N290_t2);
and AND4_12 (N485, N309_t0, N305_t0, N301_t0, N297_t0);
not NOT1_13 (N486, N405);
not NOT1_14 (N487, N44_t0);
not NOT1_15 (N488, N132_t0);
not NOT1_16 (N489, N82_t0);
not NOT1_17 (N490, N96_t0);
not NOT1_18 (N491, N69_t0);
not NOT1_19 (N492, N120_t0);
not NOT1_20 (N493, N57_t0);
not NOT1_21 (N494, N108_t0);
and AND3_22 (N495, N2_t, N15_t, N237_t0);
buf BUFF1_23 (N496, N237_t1);
and AND2_24 (N499, N37_t0, N37);
buf BUFF1_25 (N500, N219_t3);
buf BUFF1_26 (N503, N8_t0);
buf BUFF1_27 (N506, N8_t1);
buf BUFF1_28 (N509, N227_t0);
buf BUFF1_29 (N521, N234_t0);
not NOT1_30 (N533, N241_t0);
not NOT1_31 (N537, N246_t0);
and AND2_32 (N543, N11_t0, N246_t1);
and AND4_33 (N544, N132_t1, N82_t1, N96_t1, N44_t1);
and AND4_34 (N547, N120_t1, N57_t1, N108_t1, N69_t1);
buf BUFF1_35 (N550, N227_t1);
buf BUFF1_36 (N562, N234_t1);
not NOT1_37 (N574, N256_t0);
not NOT1_38 (N578, N259_t0);
buf BUFF1_39 (N582, N319_t0);
buf BUFF1_40 (N594, N322_t0);
not NOT1_41 (N606, N328_t0);
not NOT1_42 (N607, N331_t0);
not NOT1_43 (N608, N334_t0);
not NOT1_44 (N609, N337_t0);
not NOT1_45 (N610, N340_t0);
not NOT1_46 (N611, N343_t0);
not NOT1_47 (N612, N352_t0);
buf BUFF1_48 (N613, N319_t1);
buf BUFF1_49 (N625, N322_t1);
buf BUFF1_50 (N637, N16_t0);
buf BUFF1_51 (N643, N16_t1);
not NOT1_52 (N650, N355_t0);
and AND2_53 (N651, N7_t, N237_t2);
not NOT1_54 (N655, N263_t0);
not NOT1_55 (N659, N266_t0);
not NOT1_56 (N663, N269_t0);
not NOT1_57 (N667, N272_t0);
not NOT1_58 (N671, N275_t0);
not NOT1_59 (N675, N278_t0);
not NOT1_60 (N679, N281_t0);
not NOT1_61 (N683, N284_t0);
not NOT1_62 (N687, N287_t0);
buf BUFF1_63 (N693, N29_t0);
buf BUFF1_64 (N699, N29_t1);
not NOT1_65 (N705, N294_t0);
not NOT1_66 (N711, N297_t1);
not NOT1_67 (N715, N301_t1);
not NOT1_68 (N719, N305_t1);
not NOT1_69 (N723, N309_t1);
not NOT1_70 (N727, N313_t0);
not NOT1_71 (N730, N316_t0);
not NOT1_72 (N733, N346_t0);
not NOT1_73 (N734, N349_t0);
buf BUFF1_74 (N735, N259_t1);
buf BUFF1_75 (N738, N256_t1);
buf BUFF1_76 (N741, N263_t1);
buf BUFF1_77 (N744, N269_t1);
buf BUFF1_78 (N747, N266_t1);
buf BUFF1_79 (N750, N275_t1);
buf BUFF1_80 (N753, N272_t1);
buf BUFF1_81 (N756, N281_t1);
buf BUFF1_82 (N759, N278_t1);
buf BUFF1_83 (N762, N287_t1);
buf BUFF1_84 (N765, N284_t1);
buf BUFF1_85 (N768, N294_t1);
buf BUFF1_86 (N771, N301_t2);
buf BUFF1_87 (N774, N297_t2);
buf BUFF1_88 (N777, N309_t2);
buf BUFF1_89 (N780, N305_t2);
buf BUFF1_90 (N783, N316_t1);
buf BUFF1_91 (N786, N313_t1);
not NOT1_92 (N792, N485);
not NOT1_93 (N799, N495);
not NOT1_94 (N800, N499);
buf BUFF1_95 (N805, N500_t0);
nand NAND2_96 (N900, N331_t1, N606);
nand NAND2_97 (N901, N328_t1, N607);
nand NAND2_98 (N902, N337_t1, N608);
nand NAND2_99 (N903, N334_t1, N609);
nand NAND2_100 (N904, N343_t1, N610);
nand NAND2_101 (N905, N340_t1, N611);
nand NAND2_102 (N998, N349_t1, N733);
nand NAND2_103 (N999, N346_t1, N734);
and AND2_104 (N1026, N94_t, N500_t1);
and AND2_105 (N1027, N325_t0, N651_t0);
not NOT1_106 (N1028, N651_t1);
nand NAND2_107 (N1029, N231_t0, N651_t2);
not NOT1_108 (N1032, N544_t0);
not NOT1_109 (N1033, N547_t0);
and AND2_110 (N1034, N547_t1, N544_t1);
buf BUFF1_111 (N1037, N503_t0);
not NOT1_112 (N1042, N509_t0);
not NOT1_113 (N1053, N521_t0);
and AND3_114 (N1064, N80_t, N509_t1, N521_t1);
and AND3_115 (N1065, N68_t, N509_t2, N521_t2);
and AND3_116 (N1066, N79_t, N509_t3, N521_t3);
and AND3_117 (N1067, N78_t, N509_t4, N521_t4);
and AND3_118 (N1068, N77_t, N509_t5, N521_t5);
and AND2_119 (N1069, N11_t1, N537_t0);
buf BUFF1_120 (N1070, N503_t1);
not NOT1_121 (N1075, N550_t0);
not NOT1_122 (N1086, N562_t0);
and AND3_123 (N1097, N76_t, N550_t1, N562_t1);
and AND3_124 (N1098, N75_t, N550_t2, N562_t2);
and AND3_125 (N1099, N74_t, N550_t3, N562_t3);
and AND3_126 (N1100, N73_t, N550_t4, N562_t4);
and AND3_127 (N1101, N72_t, N550_t5, N562_t5);
not NOT1_128 (N1102, N582_t0);
not NOT1_129 (N1113, N594_t0);
and AND3_130 (N1124, N114_t, N582_t1, N594_t1);
and AND3_131 (N1125, N113_t, N582_t2, N594_t2);
and AND3_132 (N1126, N112_t, N582_t3, N594_t3);
and AND3_133 (N1127, N111_t, N582_t4, N594_t4);
and AND2_134 (N1128, N582_t5, N594_t5);
nand NAND2_135 (N1129, N900, N901);
nand NAND2_136 (N1133, N902, N903);
nand NAND2_137 (N1137, N904, N905);
not NOT1_138 (N1140, N741_t0);
nand NAND2_139 (N1141, N741_t1, N612);
not NOT1_140 (N1142, N744_t0);
not NOT1_141 (N1143, N747_t0);
not NOT1_142 (N1144, N750_t0);
not NOT1_143 (N1145, N753_t0);
not NOT1_144 (N1146, N613_t0);
not NOT1_145 (N1157, N625_t0);
and AND3_146 (N1168, N118_t, N613_t1, N625_t1);
and AND3_147 (N1169, N107_t, N613_t2, N625_t2);
and AND3_148 (N1170, N117_t, N613_t3, N625_t3);
and AND3_149 (N1171, N116_t, N613_t4, N625_t4);
and AND3_150 (N1172, N115_t, N613_t5, N625_t5);
not NOT1_151 (N1173, N637_t0);
not NOT1_152 (N1178, N643_t0);
not NOT1_153 (N1184, N768_t0);
nand NAND2_154 (N1185, N768_t1, N650);
not NOT1_155 (N1186, N771_t0);
not NOT1_156 (N1187, N774_t0);
not NOT1_157 (N1188, N777_t0);
not NOT1_158 (N1189, N780_t0);
buf BUFF1_159 (N1190, N506_t0);
buf BUFF1_160 (N1195, N506_t1);
not NOT1_161 (N1200, N693_t0);
not NOT1_162 (N1205, N699_t0);
not NOT1_163 (N1210, N735_t0);
not NOT1_164 (N1211, N738_t0);
not NOT1_165 (N1212, N756_t0);
not NOT1_166 (N1213, N759_t0);
not NOT1_167 (N1214, N762_t0);
not NOT1_168 (N1215, N765_t0);
nand NAND2_169 (N1216, N998, N999);
buf BUFF1_170 (N1219, N574_t0);
buf BUFF1_171 (N1222, N578_t0);
buf BUFF1_172 (N1225, N655_t0);
buf BUFF1_173 (N1228, N659_t0);
buf BUFF1_174 (N1231, N663_t0);
buf BUFF1_175 (N1234, N667_t0);
buf BUFF1_176 (N1237, N671_t0);
buf BUFF1_177 (N1240, N675_t0);
buf BUFF1_178 (N1243, N679_t0);
buf BUFF1_179 (N1246, N683_t0);
not NOT1_180 (N1249, N783_t0);
not NOT1_181 (N1250, N786_t0);
buf BUFF1_182 (N1251, N687_t0);
buf BUFF1_183 (N1254, N705_t0);
buf BUFF1_184 (N1257, N711_t0);
buf BUFF1_185 (N1260, N715_t0);
buf BUFF1_186 (N1263, N719_t0);
buf BUFF1_187 (N1266, N723_t0);
not NOT1_188 (N1269, N1027);
and AND2_189 (N1275, N325_t1, N1032);
and AND2_190 (N1276, N231_t1, N1033);
buf BUFF1_191 (N1277, N1034_t0);
or OR2_192 (N1302, N1069, N543);
nand NAND2_193 (N1351, N352_t1, N1140);
nand NAND2_194 (N1352, N747_t1, N1142);
nand NAND2_195 (N1353, N744_t1, N1143);
nand NAND2_196 (N1354, N753_t1, N1144);
nand NAND2_197 (N1355, N750_t1, N1145);
nand NAND2_198 (N1395, N355_t1, N1184);
nand NAND2_199 (N1396, N774_t1, N1186);
nand NAND2_200 (N1397, N771_t1, N1187);
nand NAND2_201 (N1398, N780_t1, N1188);
nand NAND2_202 (N1399, N777_t1, N1189);
nand NAND2_203 (N1422, N738_t1, N1210);
nand NAND2_204 (N1423, N735_t1, N1211);
nand NAND2_205 (N1424, N759_t1, N1212);
nand NAND2_206 (N1425, N756_t1, N1213);
nand NAND2_207 (N1426, N765_t1, N1214);
nand NAND2_208 (N1427, N762_t1, N1215);
nand NAND2_209 (N1440, N786_t1, N1249);
nand NAND2_210 (N1441, N783_t1, N1250);
not NOT1_211 (N1448, N1034_t1);
not NOT1_212 (N1449, N1275);
not NOT1_213 (N1450, N1276);
and AND3_214 (N1451, N93_t, N1042_t0, N1053_t0);
and AND3_215 (N1452, N55_t, N509_t6, N1053_t1);
and AND3_216 (N1453, N67_t, N1042_t1, N521_t6);
and AND3_217 (N1454, N81_t, N1042_t2, N1053_t2);
and AND3_218 (N1455, N43_t, N509_t7, N1053_t3);
and AND3_219 (N1456, N56_t, N1042_t3, N521_t7);
and AND3_220 (N1457, N92_t, N1042_t4, N1053_t4);
and AND3_221 (N1458, N54_t, N509_t8, N1053_t5);
and AND3_222 (N1459, N66_t, N1042_t5, N521_t8);
and AND3_223 (N1460, N91_t, N1042_t6, N1053_t6);
and AND3_224 (N1461, N53_t, N509_t9, N1053_t7);
and AND3_225 (N1462, N65_t, N1042_t7, N521_t9);
and AND3_226 (N1463, N90_t, N1042_t8, N1053_t8);
and AND3_227 (N1464, N52_t, N509_t10, N1053_t9);
and AND3_228 (N1465, N64_t, N1042_t9, N521_t10);
and AND3_229 (N1466, N89_t, N1075_t0, N1086_t0);
and AND3_230 (N1467, N51_t, N550_t6, N1086_t1);
and AND3_231 (N1468, N63_t, N1075_t1, N562_t6);
and AND3_232 (N1469, N88_t, N1075_t2, N1086_t2);
and AND3_233 (N1470, N50_t, N550_t7, N1086_t3);
and AND3_234 (N1471, N62_t, N1075_t3, N562_t7);
and AND3_235 (N1472, N87_t, N1075_t4, N1086_t4);
and AND3_236 (N1473, N49_t, N550_t8, N1086_t5);
and AND2_237 (N1474, N1075_t5, N562_t8);
and AND3_238 (N1475, N86_t, N1075_t6, N1086_t6);
and AND3_239 (N1476, N48_t, N550_t9, N1086_t7);
and AND3_240 (N1477, N61_t, N1075_t7, N562_t9);
and AND3_241 (N1478, N85_t, N1075_t8, N1086_t8);
and AND3_242 (N1479, N47_t, N550_t10, N1086_t9);
and AND3_243 (N1480, N60_t, N1075_t9, N562_t10);
and AND3_244 (N1481, N138_t, N1102_t0, N1113_t0);
and AND3_245 (N1482, N102_t, N582_t6, N1113_t1);
and AND3_246 (N1483, N126_t, N1102_t1, N594_t6);
and AND3_247 (N1484, N137_t, N1102_t2, N1113_t2);
and AND3_248 (N1485, N101_t, N582_t7, N1113_t3);
and AND3_249 (N1486, N125_t, N1102_t3, N594_t7);
and AND3_250 (N1487, N136_t, N1102_t4, N1113_t4);
and AND3_251 (N1488, N100_t, N582_t8, N1113_t5);
and AND3_252 (N1489, N124_t, N1102_t5, N594_t8);
and AND3_253 (N1490, N135_t, N1102_t6, N1113_t6);
and AND3_254 (N1491, N99_t, N582_t9, N1113_t7);
and AND3_255 (N1492, N123_t, N1102_t7, N594_t9);
and AND2_256 (N1493, N1102_t8, N1113_t8);
and AND2_257 (N1494, N582_t10, N1113_t9);
and AND2_258 (N1495, N1102_t9, N594_t10);
not NOT1_259 (N1496, N1129_t0);
not NOT1_260 (N1499, N1133_t0);
nand NAND2_261 (N1502, N1351, N1141);
nand NAND2_262 (N1506, N1352, N1353);
nand NAND2_263 (N1510, N1354, N1355);
buf BUFF1_264 (N1513, N1137_t0);
buf BUFF1_265 (N1516, N1137_t1);
not NOT1_266 (N1519, N1219_t0);
not NOT1_267 (N1520, N1222_t0);
not NOT1_268 (N1521, N1225_t0);
not NOT1_269 (N1522, N1228_t0);
not NOT1_270 (N1523, N1231_t0);
not NOT1_271 (N1524, N1234_t0);
not NOT1_272 (N1525, N1237_t0);
not NOT1_273 (N1526, N1240_t0);
not NOT1_274 (N1527, N1243_t0);
not NOT1_275 (N1528, N1246_t0);
and AND3_276 (N1529, N142_t, N1146_t0, N1157_t0);
and AND3_277 (N1530, N106_t, N613_t6, N1157_t1);
and AND3_278 (N1531, N130_t, N1146_t1, N625_t6);
and AND3_279 (N1532, N131_t, N1146_t2, N1157_t2);
and AND3_280 (N1533, N95_t, N613_t7, N1157_t3);
and AND3_281 (N1534, N119_t, N1146_t3, N625_t7);
and AND3_282 (N1535, N141_t, N1146_t4, N1157_t4);
and AND3_283 (N1536, N105_t, N613_t8, N1157_t5);
and AND3_284 (N1537, N129_t, N1146_t5, N625_t8);
and AND3_285 (N1538, N140_t, N1146_t6, N1157_t6);
and AND3_286 (N1539, N104_t, N613_t9, N1157_t7);
and AND3_287 (N1540, N128_t, N1146_t7, N625_t9);
and AND3_288 (N1541, N139_t, N1146_t8, N1157_t8);
and AND3_289 (N1542, N103_t, N613_t10, N1157_t9);
and AND3_290 (N1543, N127_t, N1146_t9, N625_t10);
and AND2_291 (N1544, N19_t, N1173_t0);
and AND2_292 (N1545, N4_t, N1173_t1);
and AND2_293 (N1546, N20_t, N1173_t2);
and AND2_294 (N1547, N5_t, N1173_t3);
and AND2_295 (N1548, N21_t, N1178_t0);
and AND2_296 (N1549, N22_t, N1178_t1);
and AND2_297 (N1550, N23_t, N1178_t2);
and AND2_298 (N1551, N6_t, N1178_t3);
and AND2_299 (N1552, N24_t, N1178_t4);
nand NAND2_300 (N1553, N1395, N1185);
nand NAND2_301 (N1557, N1396, N1397);
nand NAND2_302 (N1561, N1398, N1399);
and AND2_303 (N1564, N25_t, N1200_t0);
and AND2_304 (N1565, N32_t, N1200_t1);
and AND2_305 (N1566, N26_t, N1200_t2);
and AND2_306 (N1567, N33_t, N1200_t3);
and AND2_307 (N1568, N27_t, N1205_t0);
and AND2_308 (N1569, N34_t, N1205_t1);
and AND2_309 (N1570, N35_t, N1205_t2);
and AND2_310 (N1571, N28_t, N1205_t3);
not NOT1_311 (N1572, N1251_t0);
not NOT1_312 (N1573, N1254_t0);
not NOT1_313 (N1574, N1257_t0);
not NOT1_314 (N1575, N1260_t0);
not NOT1_315 (N1576, N1263_t0);
not NOT1_316 (N1577, N1266_t0);
nand NAND2_317 (N1578, N1422, N1423);
not NOT1_318 (N1581, N1216_t0);
nand NAND2_319 (N1582, N1426, N1427);
nand NAND2_320 (N1585, N1424, N1425);
nand NAND2_321 (N1588, N1440, N1441);
and AND2_322 (N1591, N1449, N1450);
or OR4_323 (N1596, N1451, N1452, N1453, N1064);
or OR4_324 (N1600, N1454, N1455, N1456, N1065);
or OR4_325 (N1606, N1457, N1458, N1459, N1066);
or OR4_326 (N1612, N1460, N1461, N1462, N1067);
or OR4_327 (N1615, N1463, N1464, N1465, N1068);
or OR4_328 (N1619, N1466, N1467, N1468, N1097);
or OR4_329 (N1624, N1469, N1470, N1471, N1098);
or OR4_330 (N1628, N1472, N1473, N1474, N1099);
or OR4_331 (N1631, N1475, N1476, N1477, N1100);
or OR4_332 (N1634, N1478, N1479, N1480, N1101);
or OR4_333 (N1637, N1481, N1482, N1483, N1124);
or OR4_334 (N1642, N1484, N1485, N1486, N1125);
or OR4_335 (N1647, N1487, N1488, N1489, N1126);
or OR4_336 (N1651, N1490, N1491, N1492, N1127);
or OR4_337 (N1656, N1493, N1494, N1495, N1128);
or OR4_338 (N1676, N1532, N1533, N1534, N1169);
or OR4_339 (N1681, N1535, N1536, N1537, N1170);
or OR4_340 (N1686, N1538, N1539, N1540, N1171);
or OR4_341 (N1690, N1541, N1542, N1543, N1172);
or OR4_342 (N1708, N1529, N1530, N1531, N1168);
buf BUFF1_343 (N1726, N1591_t0);
not NOT1_344 (N1770, N1502_t0);
not NOT1_345 (N1773, N1506_t0);
not NOT1_346 (N1776, N1513_t0);
not NOT1_347 (N1777, N1516_t0);
buf BUFF1_348 (N1778, N1510_t0);
buf BUFF1_349 (N1781, N1510_t1);
and AND3_350 (N1784, N1133_t1, N1129_t1, N1513_t1);
and AND3_351 (N1785, N1499_t0, N1496_t0, N1516_t1);
not NOT1_352 (N1795, N1553_t0);
not NOT1_353 (N1798, N1557_t0);
buf BUFF1_354 (N1801, N1561_t0);
buf BUFF1_355 (N1804, N1561_t1);
not NOT1_356 (N1807, N1588_t0);
not NOT1_357 (N1808, N1578_t0);
nand NAND2_358 (N1809, N1578_t1, N1581);
not NOT1_359 (N1810, N1582_t0);
not NOT1_360 (N1811, N1585_t0);
and AND2_361 (N1813, N1596_t0, N241_t1);
and AND2_362 (N1814, N1606_t0, N241_t2);
and AND2_363 (N1815, N1600_t0, N241_t3);
not NOT1_364 (N1816, N1642_t0);
not NOT1_365 (N1817, N1647_t0);
not NOT1_366 (N1818, N1637_t0);
not NOT1_367 (N1819, N1624_t0);
not NOT1_368 (N1820, N1619_t0);
not NOT1_369 (N1821, N1615_t0);
and AND4_370 (N1822, N496_t0, N224_t0, N36_t, N1591_t1);
and AND4_371 (N1823, N496_t1, N224_t1, N1591_t2, N486);
buf BUFF1_372 (N1824, N1596_t1);
not NOT1_373 (N1827, N1606_t1);
and AND2_374 (N1830, N1600_t1, N537_t1);
and AND2_375 (N1831, N1606_t2, N537_t2);
and AND2_376 (N1832, N1619_t1, N246_t2);
not NOT1_377 (N1833, N1596_t2);
not NOT1_378 (N1836, N1600_t2);
not NOT1_379 (N1841, N1606_t3);
buf BUFF1_380 (N1848, N1612_t0);
buf BUFF1_381 (N1852, N1615_t1);
buf BUFF1_382 (N1856, N1619_t2);
buf BUFF1_383 (N1863, N1624_t1);
buf BUFF1_384 (N1870, N1628_t0);
buf BUFF1_385 (N1875, N1631_t0);
buf BUFF1_386 (N1880, N1634_t0);
nand NAND2_387 (N1885, N727_t0, N1651_t0);
nand NAND2_388 (N1888, N730_t0, N1656_t0);
buf BUFF1_389 (N1891, N1686_t0);
and AND2_390 (N1894, N1637_t1, N425);
not NOT1_391 (N1897, N1642_t1);
and AND3_392 (N1908, N1496_t1, N1133_t2, N1776);
and AND3_393 (N1909, N1129_t2, N1499_t1, N1777);
and AND2_394 (N1910, N1600_t3, N637_t1);
and AND2_395 (N1911, N1606_t4, N637_t2);
and AND2_396 (N1912, N1612_t1, N637_t3);
and AND2_397 (N1913, N1615_t2, N637_t4);
and AND2_398 (N1914, N1619_t3, N643_t1);
and AND2_399 (N1915, N1624_t2, N643_t2);
and AND2_400 (N1916, N1628_t1, N643_t3);
and AND2_401 (N1917, N1631_t1, N643_t4);
and AND2_402 (N1918, N1634_t1, N643_t5);
not NOT1_403 (N1919, N1708_t0);
and AND2_404 (N1928, N1676_t0, N693_t1);
and AND2_405 (N1929, N1681_t0, N693_t2);
and AND2_406 (N1930, N1686_t1, N693_t3);
and AND2_407 (N1931, N1690_t0, N693_t4);
and AND2_408 (N1932, N1637_t2, N699_t1);
and AND2_409 (N1933, N1642_t2, N699_t2);
and AND2_410 (N1934, N1647_t1, N699_t3);
and AND2_411 (N1935, N1651_t1, N699_t4);
buf BUFF1_412 (N1936, N1600_t4);
nand NAND2_413 (N1939, N1216_t1, N1808);
nand NAND2_414 (N1940, N1585_t1, N1810);
nand NAND2_415 (N1941, N1582_t1, N1811);
buf BUFF1_416 (N1942, N1676_t1);
buf BUFF1_417 (N1945, N1686_t2);
buf BUFF1_418 (N1948, N1681_t1);
buf BUFF1_419 (N1951, N1637_t3);
buf BUFF1_420 (N1954, N1690_t1);
buf BUFF1_421 (N1957, N1647_t2);
buf BUFF1_422 (N1960, N1642_t3);
buf BUFF1_423 (N1963, N1656_t1);
buf BUFF1_424 (N1966, N1651_t2);
or OR2_425 (N1969, N533_t0, N1815);
not NOT1_426 (N1970, N1822);
not NOT1_427 (N1971, N1823);
buf BUFF1_428 (N2010, N1848_t0);
buf BUFF1_429 (N2012, N1852_t0);
buf BUFF1_430 (N2014, N1856_t0);
buf BUFF1_431 (N2016, N1863_t0);
buf BUFF1_432 (N2018, N1870_t0);
buf BUFF1_433 (N2020, N1875_t0);
buf BUFF1_434 (N2022, N1880_t0);
not NOT1_435 (N2028, N1778_t0);
not NOT1_436 (N2029, N1781_t0);
nor NOR2_437 (N2030, N1908, N1784);
nor NOR2_438 (N2031, N1909, N1785);
and AND3_439 (N2032, N1506_t1, N1502_t1, N1778_t1);
and AND3_440 (N2033, N1773_t0, N1770_t0, N1781_t1);
or OR2_441 (N2034, N1571, N1935);
not NOT1_442 (N2040, N1801_t0);
not NOT1_443 (N2041, N1804_t0);
and AND3_444 (N2042, N1557_t1, N1553_t1, N1801_t1);
and AND3_445 (N2043, N1798_t0, N1795_t0, N1804_t1);
nand NAND2_446 (N2046, N1939, N1809);
nand NAND2_447 (N2049, N1940, N1941);
or OR2_448 (N2052, N1544, N1910);
or OR2_449 (N2055, N1545, N1911);
or OR2_450 (N2058, N1546, N1912);
or OR2_451 (N2061, N1547, N1913);
or OR2_452 (N2064, N1548, N1914);
or OR2_453 (N2067, N1549, N1915);
or OR2_454 (N2070, N1550, N1916);
or OR2_455 (N2073, N1551, N1917);
or OR2_456 (N2076, N1552, N1918);
or OR2_457 (N2079, N1564, N1928);
or OR2_458 (N2095, N1565, N1929);
or OR2_459 (N2098, N1566, N1930);
or OR2_460 (N2101, N1567, N1931);
or OR2_461 (N2104, N1568, N1932);
or OR2_462 (N2107, N1569, N1933);
or OR2_463 (N2110, N1570, N1934);
and AND3_464 (N2113, N1897_t0, N1894_t0, N40_t0);
not NOT1_465 (N2119, N1894_t1);
nand NAND2_466 (N2120, N408, N1827_t0);
and AND2_467 (N2125, N1824_t0, N537_t3);
and AND2_468 (N2126, N1852_t1, N246_t3);
and AND2_469 (N2127, N1848_t1, N537_t4);
not NOT1_470 (N2128, N1848_t2);
not NOT1_471 (N2135, N1852_t2);
not NOT1_472 (N2141, N1863_t1);
not NOT1_473 (N2144, N1870_t1);
not NOT1_474 (N2147, N1875_t1);
not NOT1_475 (N2150, N1880_t1);
and AND2_476 (N2153, N727_t1, N1885_t0);
and AND2_477 (N2154, N1885_t1, N1651_t3);
and AND2_478 (N2155, N730_t1, N1888_t0);
and AND2_479 (N2156, N1888_t1, N1656_t2);
and AND3_480 (N2157, N1770_t1, N1506_t2, N2028);
and AND3_481 (N2158, N1502_t2, N1773_t1, N2029);
not NOT1_482 (N2171, N1942_t0);
nand NAND2_483 (N2172, N1942_t1, N1919);
not NOT1_484 (N2173, N1945_t0);
not NOT1_485 (N2174, N1948_t0);
not NOT1_486 (N2175, N1951_t0);
not NOT1_487 (N2176, N1954_t0);
and AND3_488 (N2177, N1795_t1, N1557_t2, N2040);
and AND3_489 (N2178, N1553_t2, N1798_t1, N2041);
buf BUFF1_490 (N2185, N1836_t0);
buf BUFF1_491 (N2188, N1833_t0);
buf BUFF1_492 (N2191, N1841_t0);
not NOT1_493 (N2194, N1856_t1);
not NOT1_494 (N2197, N1827_t1);
not NOT1_495 (N2200, N1936_t0);
buf BUFF1_496 (N2201, N1836_t1);
buf BUFF1_497 (N2204, N1833_t1);
buf BUFF1_498 (N2207, N1841_t1);
buf BUFF1_499 (N2210, N1824_t1);
buf BUFF1_500 (N2213, N1841_t2);
buf BUFF1_501 (N2216, N1841_t3);
nand NAND2_502 (N2219, N2031, N2030);
not NOT1_503 (N2234, N1957_t0);
not NOT1_504 (N2235, N1960_t0);
not NOT1_505 (N2236, N1963_t0);
not NOT1_506 (N2237, N1966_t0);
and AND3_507 (N2250, N40_t1, N1897_t1, N2119);
or OR2_508 (N2266, N1831, N2126);
or OR2_509 (N2269, N2127, N1832);
or OR2_510 (N2291, N2153, N2154);
or OR2_511 (N2294, N2155, N2156);
nor NOR2_512 (N2297, N2157, N2032);
nor NOR2_513 (N2298, N2158, N2033);
not NOT1_514 (N2300, N2046_t0);
not NOT1_515 (N2301, N2049_t0);
nand NAND2_516 (N2302, N2052_t0, N1519);
not NOT1_517 (N2303, N2052_t1);
nand NAND2_518 (N2304, N2055_t0, N1520);
not NOT1_519 (N2305, N2055_t1);
nand NAND2_520 (N2306, N2058_t0, N1521);
not NOT1_521 (N2307, N2058_t1);
nand NAND2_522 (N2308, N2061_t0, N1522);
not NOT1_523 (N2309, N2061_t1);
nand NAND2_524 (N2310, N2064_t0, N1523);
not NOT1_525 (N2311, N2064_t1);
nand NAND2_526 (N2312, N2067_t0, N1524);
not NOT1_527 (N2313, N2067_t1);
nand NAND2_528 (N2314, N2070_t0, N1525);
not NOT1_529 (N2315, N2070_t1);
nand NAND2_530 (N2316, N2073_t0, N1526);
not NOT1_531 (N2317, N2073_t1);
nand NAND2_532 (N2318, N2076_t0, N1527);
not NOT1_533 (N2319, N2076_t1);
nand NAND2_534 (N2320, N2079_t0, N1528);
not NOT1_535 (N2321, N2079_t1);
nand NAND2_536 (N2322, N1708_t1, N2171);
nand NAND2_537 (N2323, N1948_t1, N2173);
nand NAND2_538 (N2324, N1945_t1, N2174);
nand NAND2_539 (N2325, N1954_t1, N2175);
nand NAND2_540 (N2326, N1951_t1, N2176);
nor NOR2_541 (N2327, N2177, N2042);
nor NOR2_542 (N2328, N2178, N2043);
nand NAND2_543 (N2329, N2095_t0, N1572);
not NOT1_544 (N2330, N2095_t1);
nand NAND2_545 (N2331, N2098_t0, N1573);
not NOT1_546 (N2332, N2098_t1);
nand NAND2_547 (N2333, N2101_t0, N1574);
not NOT1_548 (N2334, N2101_t1);
nand NAND2_549 (N2335, N2104_t0, N1575);
not NOT1_550 (N2336, N2104_t1);
nand NAND2_551 (N2337, N2107_t0, N1576);
not NOT1_552 (N2338, N2107_t1);
nand NAND2_553 (N2339, N2110_t0, N1577);
not NOT1_554 (N2340, N2110_t1);
nand NAND2_555 (N2354, N1960_t1, N2234);
nand NAND2_556 (N2355, N1957_t1, N2235);
nand NAND2_557 (N2356, N1966_t1, N2236);
nand NAND2_558 (N2357, N1963_t1, N2237);
and AND2_559 (N2358, N2120_t0, N533_t1);
not NOT1_560 (N2359, N2113_t0);
not NOT1_561 (N2364, N2185_t0);
not NOT1_562 (N2365, N2188_t0);
not NOT1_563 (N2366, N2191_t0);
not NOT1_564 (N2367, N2194_t0);
buf BUFF1_565 (N2368, N2120_t1);
not NOT1_566 (N2372, N2201_t0);
not NOT1_567 (N2373, N2204_t0);
not NOT1_568 (N2374, N2207_t0);
not NOT1_569 (N2375, N2210_t0);
not NOT1_570 (N2376, N2213_t0);
not NOT1_571 (N2377, N2113_t1);
buf BUFF1_572 (N2382, N2113_t2);
and AND2_573 (N2386, N2120_t2, N246_t4);
buf BUFF1_574 (N2387, N2266_t0);
buf BUFF1_575 (N2388, N2266_t1);
buf BUFF1_576 (N2389, N2269_t0);
buf BUFF1_577 (N2390, N2269_t1);
buf BUFF1_578 (N2391, N2113_t3);
not NOT1_579 (N2395, N2113_t4);
nand NAND2_580 (N2400, N2219_t0, N2300);
not NOT1_581 (N2403, N2216_t0);
not NOT1_582 (N2406, N2219_t1);
nand NAND2_583 (N2407, N1219_t1, N2303);
nand NAND2_584 (N2408, N1222_t1, N2305);
nand NAND2_585 (N2409, N1225_t1, N2307);
nand NAND2_586 (N2410, N1228_t1, N2309);
nand NAND2_587 (N2411, N1231_t1, N2311);
nand NAND2_588 (N2412, N1234_t1, N2313);
nand NAND2_589 (N2413, N1237_t1, N2315);
nand NAND2_590 (N2414, N1240_t1, N2317);
nand NAND2_591 (N2415, N1243_t1, N2319);
nand NAND2_592 (N2416, N1246_t1, N2321);
nand NAND2_593 (N2417, N2322, N2172);
nand NAND2_594 (N2421, N2323, N2324);
nand NAND2_595 (N2425, N2325, N2326);
nand NAND2_596 (N2428, N1251_t1, N2330);
nand NAND2_597 (N2429, N1254_t1, N2332);
nand NAND2_598 (N2430, N1257_t1, N2334);
nand NAND2_599 (N2431, N1260_t1, N2336);
nand NAND2_600 (N2432, N1263_t1, N2338);
nand NAND2_601 (N2433, N1266_t1, N2340);
buf BUFF1_602 (N2434, N2128_t0);
buf BUFF1_603 (N2437, N2135_t0);
buf BUFF1_604 (N2440, N2144_t0);
buf BUFF1_605 (N2443, N2141_t0);
buf BUFF1_606 (N2446, N2150_t0);
buf BUFF1_607 (N2449, N2147_t0);
not NOT1_608 (N2452, N2197_t0);
nand NAND2_609 (N2453, N2197_t1, N2200);
buf BUFF1_610 (N2454, N2128_t1);
buf BUFF1_611 (N2457, N2144_t1);
buf BUFF1_612 (N2460, N2141_t1);
buf BUFF1_613 (N2463, N2150_t1);
buf BUFF1_614 (N2466, N2147_t1);
not NOT1_615 (N2469, N2120_t3);
buf BUFF1_616 (N2472, N2128_t2);
buf BUFF1_617 (N2475, N2135_t1);
buf BUFF1_618 (N2478, N2128_t3);
buf BUFF1_619 (N2481, N2135_t2);
nand NAND2_620 (N2484, N2298, N2297);
nand NAND2_621 (N2487, N2356, N2357);
nand NAND2_622 (N2490, N2354, N2355);
nand NAND2_623 (N2493, N2328, N2327);
or OR2_624 (N2496, N2358, N1814);
nand NAND2_625 (N2503, N2188_t1, N2364);
nand NAND2_626 (N2504, N2185_t1, N2365);
nand NAND2_627 (N2510, N2204_t1, N2372);
nand NAND2_628 (N2511, N2201_t1, N2373);
or OR2_629 (N2521, N1830, N2386);
nand NAND2_630 (N2528, N2046_t1, N2406);
not NOT1_631 (N2531, N2291_t0);
not NOT1_632 (N2534, N2294_t0);
buf BUFF1_633 (N2537, N2250_t0);
buf BUFF1_634 (N2540, N2250_t1);
nand NAND2_635 (N2544, N2302, N2407);
nand NAND2_636 (N2545, N2304, N2408);
nand NAND2_637 (N2546, N2306, N2409);
nand NAND2_638 (N2547, N2308, N2410);
nand NAND2_639 (N2548, N2310, N2411);
nand NAND2_640 (N2549, N2312, N2412);
nand NAND2_641 (N2550, N2314, N2413);
nand NAND2_642 (N2551, N2316, N2414);
nand NAND2_643 (N2552, N2318, N2415);
nand NAND2_644 (N2553, N2320, N2416);
nand NAND2_645 (N2563, N2329, N2428);
nand NAND2_646 (N2564, N2331, N2429);
nand NAND2_647 (N2565, N2333, N2430);
nand NAND2_648 (N2566, N2335, N2431);
nand NAND2_649 (N2567, N2337, N2432);
nand NAND2_650 (N2568, N2339, N2433);
nand NAND2_651 (N2579, N1936_t1, N2452);
buf BUFF1_652 (N2603, N2359_t0);
and AND2_653 (N2607, N1880_t2, N2377_t0);
and AND2_654 (N2608, N1676_t2, N2377_t1);
and AND2_655 (N2609, N1681_t2, N2377_t2);
and AND2_656 (N2610, N1891_t0, N2377_t3);
and AND2_657 (N2611, N1856_t2, N2382_t0);
and AND2_658 (N2612, N1863_t2, N2382_t1);
nand NAND2_659 (N2613, N2503, N2504);
not NOT1_660 (N2617, N2434_t0);
nand NAND2_661 (N2618, N2434_t1, N2366);
nand NAND2_662 (N2619, N2437_t0, N2367);
not NOT1_663 (N2620, N2437_t1);
not NOT1_664 (N2621, N2368_t0);
nand NAND2_665 (N2624, N2510, N2511);
not NOT1_666 (N2628, N2454_t0);
nand NAND2_667 (N2629, N2454_t1, N2374);
not NOT1_668 (N2630, N2472_t0);
and AND2_669 (N2631, N1856_t3, N2391_t0);
and AND2_670 (N2632, N1863_t3, N2391_t1);
and AND2_671 (N2633, N1880_t3, N2395_t0);
and AND2_672 (N2634, N1676_t3, N2395_t1);
and AND2_673 (N2635, N1681_t3, N2395_t2);
and AND2_674 (N2636, N1891_t1, N2395_t3);
not NOT1_675 (N2638, N2382_t2);
buf BUFF1_676 (N2643, N2521_t0);
buf BUFF1_677 (N2644, N2521_t1);
not NOT1_678 (N2645, N2475_t0);
not NOT1_679 (N2646, N2391_t2);
nand NAND2_680 (N2652, N2528, N2400);
not NOT1_681 (N2655, N2478_t0);
not NOT1_682 (N2656, N2481_t0);
buf BUFF1_683 (N2659, N2359_t1);
not NOT1_684 (N2663, N2484_t0);
nand NAND2_685 (N2664, N2484_t1, N2301);
not NOT1_686 (N2665, N2553);
not NOT1_687 (N2666, N2552);
not NOT1_688 (N2667, N2551);
not NOT1_689 (N2668, N2550);
not NOT1_690 (N2669, N2549);
not NOT1_691 (N2670, N2548);
not NOT1_692 (N2671, N2547);
not NOT1_693 (N2672, N2546);
not NOT1_694 (N2673, N2545);
not NOT1_695 (N2674, N2544);
not NOT1_696 (N2675, N2568);
not NOT1_697 (N2676, N2567);
not NOT1_698 (N2677, N2566);
not NOT1_699 (N2678, N2565);
not NOT1_700 (N2679, N2564);
not NOT1_701 (N2680, N2563);
not NOT1_702 (N2681, N2417_t0);
not NOT1_703 (N2684, N2421_t0);
buf BUFF1_704 (N2687, N2425_t0);
buf BUFF1_705 (N2690, N2425_t1);
not NOT1_706 (N2693, N2493_t0);
nand NAND2_707 (N2694, N2493_t1, N1807);
not NOT1_708 (N2695, N2440_t0);
not NOT1_709 (N2696, N2443_t0);
not NOT1_710 (N2697, N2446_t0);
not NOT1_711 (N2698, N2449_t0);
not NOT1_712 (N2699, N2457_t0);
not NOT1_713 (N2700, N2460_t0);
not NOT1_714 (N2701, N2463_t0);
not NOT1_715 (N2702, N2466_t0);
nand NAND2_716 (N2703, N2579, N2453);
not NOT1_717 (N2706, N2469_t0);
not NOT1_718 (N2707, N2487_t0);
not NOT1_719 (N2708, N2490_t0);
and AND2_720 (N2709, N2294_t1, N2534_t0);
and AND2_721 (N2710, N2291_t1, N2531_t0);
nand NAND2_722 (N2719, N2191_t1, N2617);
nand NAND2_723 (N2720, N2194_t1, N2620);
nand NAND2_724 (N2726, N2207_t1, N2628);
buf BUFF1_725 (N2729, N2537_t0);
buf BUFF1_726 (N2738, N2537_t1);
not NOT1_727 (N2743, N2652);
nand NAND2_728 (N2747, N2049_t1, N2663);
and AND5_729 (N2748, N2665, N2666, N2667, N2668, N2669);
and AND5_730 (N2749, N2670, N2671, N2672, N2673, N2674);
and AND2_731 (N2750, N2034, N2675);
and AND5_732 (N2751, N2676, N2677, N2678, N2679, N2680);
nand NAND2_733 (N2760, N1588_t1, N2693);
buf BUFF1_734 (N2761, N2540_t0);
buf BUFF1_735 (N2766, N2540_t1);
nand NAND2_736 (N2771, N2443_t1, N2695);
nand NAND2_737 (N2772, N2440_t1, N2696);
nand NAND2_738 (N2773, N2449_t1, N2697);
nand NAND2_739 (N2774, N2446_t1, N2698);
nand NAND2_740 (N2775, N2460_t1, N2699);
nand NAND2_741 (N2776, N2457_t1, N2700);
nand NAND2_742 (N2777, N2466_t1, N2701);
nand NAND2_743 (N2778, N2463_t1, N2702);
nand NAND2_744 (N2781, N2490_t1, N2707);
nand NAND2_745 (N2782, N2487_t1, N2708);
or OR2_746 (N2783, N2709, N2534_t1);
or OR2_747 (N2784, N2710, N2531_t1);
and AND2_748 (N2789, N1856_t4, N2638_t0);
and AND2_749 (N2790, N1863_t4, N2638_t1);
and AND2_750 (N2791, N1870_t2, N2638_t2);
and AND2_751 (N2792, N1875_t2, N2638_t3);
not NOT1_752 (N2793, N2613_t0);
nand NAND2_753 (N2796, N2719, N2618);
nand NAND2_754 (N2800, N2619, N2720);
not NOT1_755 (N2803, N2624_t0);
nand NAND2_756 (N2806, N2726, N2629);
and AND2_757 (N2809, N1856_t5, N2646_t0);
and AND2_758 (N2810, N1863_t5, N2646_t1);
and AND2_759 (N2811, N1870_t3, N2646_t2);
and AND2_760 (N2812, N1875_t3, N2646_t3);
and AND2_761 (N2817, N2743, N14_t);
buf BUFF1_762 (N2820, N2603_t0);
nand NAND2_763 (N2826, N2747, N2664);
and AND2_764 (N2829, N2748, N2749);
and AND2_765 (N2830, N2750, N2751);
buf BUFF1_766 (N2831, N2659_t0);
not NOT1_767 (N2837, N2687_t0);
not NOT1_768 (N2838, N2690_t0);
and AND3_769 (N2839, N2421_t1, N2417_t1, N2687_t1);
and AND3_770 (N2840, N2684_t0, N2681_t0, N2690_t1);
nand NAND2_771 (N2841, N2760, N2694);
buf BUFF1_772 (N2844, N2603_t1);
buf BUFF1_773 (N2854, N2603_t2);
buf BUFF1_774 (N2859, N2659_t1);
buf BUFF1_775 (N2869, N2659_t2);
nand NAND2_776 (N2874, N2773, N2774);
nand NAND2_777 (N2877, N2771, N2772);
not NOT1_778 (N2880, N2703_t0);
nand NAND2_779 (N2881, N2703_t1, N2706);
nand NAND2_780 (N2882, N2777, N2778);
nand NAND2_781 (N2885, N2775, N2776);
nand NAND2_782 (N2888, N2781, N2782);
nand NAND2_783 (N2891, N2783, N2784);
and AND2_784 (N2894, N2607, N2729_t0);
and AND2_785 (N2895, N2608, N2729_t1);
and AND2_786 (N2896, N2609, N2729_t2);
and AND2_787 (N2897, N2610, N2729_t3);
or OR2_788 (N2898, N2789, N2611);
or OR2_789 (N2899, N2790, N2612);
and AND2_790 (N2900, N2791, N1037_t0);
and AND2_791 (N2901, N2792, N1037_t1);
or OR2_792 (N2914, N2809, N2631);
or OR2_793 (N2915, N2810, N2632);
and AND2_794 (N2916, N2811, N1070_t0);
and AND2_795 (N2917, N2812, N1070_t1);
and AND2_796 (N2918, N2633, N2738_t0);
and AND2_797 (N2919, N2634, N2738_t1);
and AND2_798 (N2920, N2635, N2738_t2);
and AND2_799 (N2921, N2636, N2738_t3);
buf BUFF1_800 (N2925, N2817_t0);
and AND3_801 (N2931, N2829, N2830, N1302);
and AND3_802 (N2938, N2681_t1, N2421_t2, N2837);
and AND3_803 (N2939, N2417_t2, N2684_t1, N2838);
nand NAND2_804 (N2963, N2469_t1, N2880);
not NOT1_805 (N2970, N2841_t0);
not NOT1_806 (N2971, N2826_t0);
not NOT1_807 (N2972, N2894);
not NOT1_808 (N2975, N2895);
not NOT1_809 (N2978, N2896);
not NOT1_810 (N2981, N2897);
and AND2_811 (N2984, N2898, N1037_t2);
and AND2_812 (N2985, N2899, N1037_t3);
not NOT1_813 (N2986, N2900);
not NOT1_814 (N2989, N2901);
not NOT1_815 (N2992, N2796_t0);
buf BUFF1_816 (N2995, N2800_t0);
buf BUFF1_817 (N2998, N2800_t1);
buf BUFF1_818 (N3001, N2806_t0);
buf BUFF1_819 (N3004, N2806_t1);
and AND2_820 (N3007, N574_t1, N2820_t0);
and AND2_821 (N3008, N2914, N1070_t2);
and AND2_822 (N3009, N2915, N1070_t3);
not NOT1_823 (N3010, N2916);
not NOT1_824 (N3013, N2917);
not NOT1_825 (N3016, N2918);
not NOT1_826 (N3019, N2919);
not NOT1_827 (N3022, N2920);
not NOT1_828 (N3025, N2921);
not NOT1_829 (N3028, N2817_t1);
and AND2_830 (N3029, N574_t2, N2831_t0);
not NOT1_831 (N3030, N2820_t1);
and AND2_832 (N3035, N578_t1, N2820_t2);
and AND2_833 (N3036, N655_t1, N2820_t3);
and AND2_834 (N3037, N659_t1, N2820_t4);
buf BUFF1_835 (N3038, N2931_t0);
not NOT1_836 (N3039, N2831_t1);
and AND2_837 (N3044, N578_t2, N2831_t2);
and AND2_838 (N3045, N655_t2, N2831_t3);
and AND2_839 (N3046, N659_t2, N2831_t4);
nor NOR2_840 (N3047, N2938, N2839);
nor NOR2_841 (N3048, N2939, N2840);
not NOT1_842 (N3049, N2888_t0);
not NOT1_843 (N3050, N2844_t0);
and AND2_844 (N3053, N663_t1, N2844_t1);
and AND2_845 (N3054, N667_t1, N2844_t2);
and AND2_846 (N3055, N671_t1, N2844_t3);
and AND2_847 (N3056, N675_t1, N2844_t4);
and AND2_848 (N3057, N679_t1, N2854_t0);
and AND2_849 (N3058, N683_t1, N2854_t1);
and AND2_850 (N3059, N687_t1, N2854_t2);
and AND2_851 (N3060, N705_t1, N2854_t3);
not NOT1_852 (N3061, N2859_t0);
and AND2_853 (N3064, N663_t2, N2859_t1);
and AND2_854 (N3065, N667_t2, N2859_t2);
and AND2_855 (N3066, N671_t2, N2859_t3);
and AND2_856 (N3067, N675_t2, N2859_t4);
and AND2_857 (N3068, N679_t2, N2869_t0);
and AND2_858 (N3069, N683_t2, N2869_t1);
and AND2_859 (N3070, N687_t2, N2869_t2);
and AND2_860 (N3071, N705_t2, N2869_t3);
not NOT1_861 (N3072, N2874_t0);
not NOT1_862 (N3073, N2877_t0);
not NOT1_863 (N3074, N2882_t0);
not NOT1_864 (N3075, N2885_t0);
nand NAND2_865 (N3076, N2881, N2963);
not NOT1_866 (N3079, N2931_t1);
not NOT1_867 (N3088, N2984);
not NOT1_868 (N3091, N2985);
not NOT1_869 (N3110, N3008);
not NOT1_870 (N3113, N3009);
and AND2_871 (N3137, N3055, N1190_t0);
and AND2_872 (N3140, N3056, N1190_t1);
and AND2_873 (N3143, N3057, N2761_t0);
and AND2_874 (N3146, N3058, N2761_t1);
and AND2_875 (N3149, N3059, N2761_t2);
and AND2_876 (N3152, N3060, N2761_t3);
and AND2_877 (N3157, N3066, N1195_t0);
and AND2_878 (N3160, N3067, N1195_t1);
and AND2_879 (N3163, N3068, N2766_t0);
and AND2_880 (N3166, N3069, N2766_t1);
and AND2_881 (N3169, N3070, N2766_t2);
and AND2_882 (N3172, N3071, N2766_t3);
nand NAND2_883 (N3175, N2877_t1, N3072);
nand NAND2_884 (N3176, N2874_t1, N3073);
nand NAND2_885 (N3177, N2885_t1, N3074);
nand NAND2_886 (N3178, N2882_t1, N3075);
nand NAND2_887 (N3180, N3048, N3047);
not NOT1_888 (N3187, N2995_t0);
not NOT1_889 (N3188, N2998_t0);
not NOT1_890 (N3189, N3001_t0);
not NOT1_891 (N3190, N3004_t0);
and AND3_892 (N3191, N2796_t1, N2613_t1, N2995_t1);
and AND3_893 (N3192, N2992_t0, N2793_t0, N2998_t1);
and AND3_894 (N3193, N2624_t1, N2368_t1, N3001_t1);
and AND3_895 (N3194, N2803_t0, N2621_t0, N3004_t1);
nand NAND2_896 (N3195, N3076_t0, N2375);
not NOT1_897 (N3196, N3076_t1);
and AND2_898 (N3197, N687_t3, N3030_t0);
and AND2_899 (N3208, N687_t4, N3039_t0);
and AND2_900 (N3215, N705_t3, N3030_t1);
and AND2_901 (N3216, N711_t1, N3030_t2);
and AND2_902 (N3217, N715_t1, N3030_t3);
and AND2_903 (N3218, N705_t4, N3039_t1);
and AND2_904 (N3219, N711_t2, N3039_t2);
and AND2_905 (N3220, N715_t2, N3039_t3);
and AND2_906 (N3222, N719_t1, N3050_t0);
and AND2_907 (N3223, N723_t1, N3050_t1);
and AND2_908 (N3230, N719_t2, N3061_t0);
and AND2_909 (N3231, N723_t2, N3061_t1);
nand NAND2_910 (N3238, N3175, N3176);
nand NAND2_911 (N3241, N3177, N3178);
buf BUFF1_912 (N3244, N2981_t0);
buf BUFF1_913 (N3247, N2978_t0);
buf BUFF1_914 (N3250, N2975_t0);
buf BUFF1_915 (N3253, N2972_t0);
buf BUFF1_916 (N3256, N2989_t0);
buf BUFF1_917 (N3259, N2986_t0);
buf BUFF1_918 (N3262, N3025_t0);
buf BUFF1_919 (N3265, N3022_t0);
buf BUFF1_920 (N3268, N3019_t0);
buf BUFF1_921 (N3271, N3016_t0);
buf BUFF1_922 (N3274, N3013_t0);
buf BUFF1_923 (N3277, N3010_t0);
and AND3_924 (N3281, N2793_t1, N2796_t2, N3187);
and AND3_925 (N3282, N2613_t2, N2992_t1, N3188);
and AND3_926 (N3283, N2621_t1, N2624_t2, N3189);
and AND3_927 (N3284, N2368_t2, N2803_t1, N3190);
nand NAND2_928 (N3286, N2210_t1, N3196);
or OR2_929 (N3288, N3197, N3007);
nand NAND2_930 (N3289, N3180_t0, N3049);
and AND2_931 (N3291, N3152_t0, N2981_t1);
and AND2_932 (N3293, N3149_t0, N2978_t1);
and AND2_933 (N3295, N3146_t0, N2975_t1);
and AND2_934 (N3296, N2972_t1, N3143_t0);
and AND2_935 (N3299, N3140_t0, N2989_t1);
and AND2_936 (N3301, N3137_t0, N2986_t1);
or OR2_937 (N3302, N3208, N3029);
and AND2_938 (N3304, N3172_t0, N3025_t1);
and AND2_939 (N3306, N3169_t0, N3022_t1);
and AND2_940 (N3308, N3166_t0, N3019_t1);
and AND2_941 (N3309, N3016_t1, N3163_t0);
and AND2_942 (N3312, N3160_t0, N3013_t1);
and AND2_943 (N3314, N3157_t0, N3010_t1);
or OR2_944 (N3315, N3215, N3035);
or OR2_945 (N3318, N3216, N3036);
or OR2_946 (N3321, N3217, N3037);
or OR2_947 (N3324, N3218, N3044);
or OR2_948 (N3327, N3219, N3045);
or OR2_949 (N3330, N3220, N3046);
not NOT1_950 (N3333, N3180_t1);
or OR2_951 (N3334, N3222, N3053);
or OR2_952 (N3335, N3223, N3054);
or OR2_953 (N3336, N3230, N3064);
or OR2_954 (N3337, N3231, N3065);
buf BUFF1_955 (N3340, N3152_t1);
buf BUFF1_956 (N3344, N3149_t1);
buf BUFF1_957 (N3348, N3146_t1);
buf BUFF1_958 (N3352, N3143_t1);
buf BUFF1_959 (N3356, N3140_t1);
buf BUFF1_960 (N3360, N3137_t1);
buf BUFF1_961 (N3364, N3091_t0);
buf BUFF1_962 (N3367, N3088_t0);
buf BUFF1_963 (N3370, N3172_t1);
buf BUFF1_964 (N3374, N3169_t1);
buf BUFF1_965 (N3378, N3166_t1);
buf BUFF1_966 (N3382, N3163_t1);
buf BUFF1_967 (N3386, N3160_t1);
buf BUFF1_968 (N3390, N3157_t1);
buf BUFF1_969 (N3394, N3113_t0);
buf BUFF1_970 (N3397, N3110_t0);
nand NAND2_971 (N3400, N3195, N3286);
nor NOR2_972 (N3401, N3281, N3191);
nor NOR2_973 (N3402, N3282, N3192);
nor NOR2_974 (N3403, N3283, N3193);
nor NOR2_975 (N3404, N3284, N3194);
not NOT1_976 (N3405, N3238_t0);
not NOT1_977 (N3406, N3241_t0);
and AND2_978 (N3409, N3288, N1836_t2);
nand NAND2_979 (N3410, N2888_t1, N3333);
not NOT1_980 (N3412, N3244_t0);
not NOT1_981 (N3414, N3247_t0);
not NOT1_982 (N3416, N3250_t0);
not NOT1_983 (N3418, N3253_t0);
not NOT1_984 (N3420, N3256_t0);
not NOT1_985 (N3422, N3259_t0);
and AND2_986 (N3428, N3302, N1836_t3);
not NOT1_987 (N3430, N3262_t0);
not NOT1_988 (N3432, N3265_t0);
not NOT1_989 (N3434, N3268_t0);
not NOT1_990 (N3436, N3271_t0);
not NOT1_991 (N3438, N3274_t0);
not NOT1_992 (N3440, N3277_t0);
and AND2_993 (N3450, N3334, N1190_t2);
and AND2_994 (N3453, N3335, N1190_t3);
and AND2_995 (N3456, N3336, N1195_t2);
and AND2_996 (N3459, N3337, N1195_t3);
and AND2_997 (N3478, N3400, N533_t2);
and AND2_998 (N3479, N3318_t0, N2128_t4);
and AND2_999 (N3480, N3315_t0, N1841_t4);
nand NAND2_1000 (N3481, N3410, N3289);
not NOT1_1001 (N3482, N3340_t0);
nand NAND2_1002 (N3483, N3340_t1, N3412);
not NOT1_1003 (N3484, N3344_t0);
nand NAND2_1004 (N3485, N3344_t1, N3414);
not NOT1_1005 (N3486, N3348_t0);
nand NAND2_1006 (N3487, N3348_t1, N3416);
not NOT1_1007 (N3488, N3352_t0);
nand NAND2_1008 (N3489, N3352_t1, N3418);
not NOT1_1009 (N3490, N3356_t0);
nand NAND2_1010 (N3491, N3356_t1, N3420);
not NOT1_1011 (N3492, N3360_t0);
nand NAND2_1012 (N3493, N3360_t1, N3422);
not NOT1_1013 (N3494, N3364_t0);
not NOT1_1014 (N3496, N3367_t0);
and AND2_1015 (N3498, N3321_t0, N2135_t3);
and AND2_1016 (N3499, N3327_t0, N2128_t5);
and AND2_1017 (N3500, N3324_t0, N1841_t5);
not NOT1_1018 (N3501, N3370_t0);
nand NAND2_1019 (N3502, N3370_t1, N3430);
not NOT1_1020 (N3503, N3374_t0);
nand NAND2_1021 (N3504, N3374_t1, N3432);
not NOT1_1022 (N3505, N3378_t0);
nand NAND2_1023 (N3506, N3378_t1, N3434);
not NOT1_1024 (N3507, N3382_t0);
nand NAND2_1025 (N3508, N3382_t1, N3436);
not NOT1_1026 (N3509, N3386_t0);
nand NAND2_1027 (N3510, N3386_t1, N3438);
not NOT1_1028 (N3511, N3390_t0);
nand NAND2_1029 (N3512, N3390_t1, N3440);
not NOT1_1030 (N3513, N3394_t0);
not NOT1_1031 (N3515, N3397_t0);
and AND2_1032 (N3517, N3330_t0, N2135_t4);
nand NAND2_1033 (N3522, N3402, N3401);
nand NAND2_1034 (N3525, N3404, N3403);
buf BUFF1_1035 (N3528, N3318_t1);
buf BUFF1_1036 (N3531, N3315_t1);
buf BUFF1_1037 (N3534, N3321_t1);
buf BUFF1_1038 (N3537, N3327_t1);
buf BUFF1_1039 (N3540, N3324_t1);
buf BUFF1_1040 (N3543, N3330_t1);
or OR2_1041 (N3546, N3478, N1813);
not NOT1_1042 (N3551, N3481);
nand NAND2_1043 (N3552, N3244_t1, N3482);
nand NAND2_1044 (N3553, N3247_t1, N3484);
nand NAND2_1045 (N3554, N3250_t1, N3486);
nand NAND2_1046 (N3555, N3253_t1, N3488);
nand NAND2_1047 (N3556, N3256_t1, N3490);
nand NAND2_1048 (N3557, N3259_t1, N3492);
and AND2_1049 (N3558, N3453_t0, N3091_t1);
and AND2_1050 (N3559, N3450_t0, N3088_t1);
nand NAND2_1051 (N3563, N3262_t1, N3501);
nand NAND2_1052 (N3564, N3265_t1, N3503);
nand NAND2_1053 (N3565, N3268_t1, N3505);
nand NAND2_1054 (N3566, N3271_t1, N3507);
nand NAND2_1055 (N3567, N3274_t1, N3509);
nand NAND2_1056 (N3568, N3277_t1, N3511);
and AND2_1057 (N3569, N3459_t0, N3113_t1);
and AND2_1058 (N3570, N3456_t0, N3110_t1);
buf BUFF1_1059 (N3576, N3453_t1);
buf BUFF1_1060 (N3579, N3450_t1);
buf BUFF1_1061 (N3585, N3459_t1);
buf BUFF1_1062 (N3588, N3456_t1);
not NOT1_1063 (N3592, N3522_t0);
nand NAND2_1064 (N3593, N3522_t1, N3405);
not NOT1_1065 (N3594, N3525_t0);
nand NAND2_1066 (N3595, N3525_t1, N3406);
not NOT1_1067 (N3596, N3528_t0);
nand NAND2_1068 (N3597, N3528_t1, N2630);
nand NAND2_1069 (N3598, N3531_t0, N2376);
not NOT1_1070 (N3599, N3531_t1);
and AND2_1071 (N3600, N3551, N800_t0);
nand NAND2_1072 (N3603, N3552, N3483);
nand NAND2_1073 (N3608, N3553, N3485);
nand NAND2_1074 (N3612, N3554, N3487);
nand NAND2_1075 (N3615, N3555, N3489);
nand NAND2_1076 (N3616, N3556, N3491);
nand NAND2_1077 (N3622, N3557, N3493);
not NOT1_1078 (N3629, N3534_t0);
nand NAND2_1079 (N3630, N3534_t1, N2645);
not NOT1_1080 (N3631, N3537_t0);
nand NAND2_1081 (N3632, N3537_t1, N2655);
nand NAND2_1082 (N3633, N3540_t0, N2403);
not NOT1_1083 (N3634, N3540_t1);
nand NAND2_1084 (N3635, N3563, N3502);
nand NAND2_1085 (N3640, N3564, N3504);
nand NAND2_1086 (N3644, N3565, N3506);
nand NAND2_1087 (N3647, N3566, N3508);
nand NAND2_1088 (N3648, N3567, N3510);
nand NAND2_1089 (N3654, N3568, N3512);
not NOT1_1090 (N3661, N3543_t0);
nand NAND2_1091 (N3662, N3543_t1, N2656);
nand NAND2_1092 (N3667, N3238_t1, N3592);
nand NAND2_1093 (N3668, N3241_t1, N3594);
nand NAND2_1094 (N3669, N2472_t1, N3596);
nand NAND2_1095 (N3670, N2213_t1, N3599);
buf BUFF1_1096 (N3671, N3600_t0);
not NOT1_1097 (N3691, N3576_t0);
nand NAND2_1098 (N3692, N3576_t1, N3494);
not NOT1_1099 (N3693, N3579_t0);
nand NAND2_1100 (N3694, N3579_t1, N3496);
nand NAND2_1101 (N3695, N2475_t1, N3629);
nand NAND2_1102 (N3696, N2478_t1, N3631);
nand NAND2_1103 (N3697, N2216_t1, N3634);
not NOT1_1104 (N3716, N3585_t0);
nand NAND2_1105 (N3717, N3585_t1, N3513);
not NOT1_1106 (N3718, N3588_t0);
nand NAND2_1107 (N3719, N3588_t1, N3515);
nand NAND2_1108 (N3720, N2481_t1, N3661);
nand NAND2_1109 (N3721, N3667, N3593);
nand NAND2_1110 (N3722, N3668, N3595);
nand NAND2_1111 (N3723, N3669, N3597);
nand NAND2_1112 (N3726, N3670, N3598);
not NOT1_1113 (N3727, N3600_t1);
nand NAND2_1114 (N3728, N3364_t1, N3691);
nand NAND2_1115 (N3729, N3367_t1, N3693);
nand NAND2_1116 (N3730, N3695, N3630);
and AND4_1117 (N3731, N3608_t0, N3615, N3612_t0, N3603_t0);
and AND2_1118 (N3732, N3603_t1, N3293);
and AND3_1119 (N3733, N3608_t1, N3603_t2, N3295);
and AND4_1120 (N3734, N3612_t1, N3603_t3, N3296, N3608_t2);
and AND2_1121 (N3735, N3616_t0, N3301);
and AND3_1122 (N3736, N3622_t0, N3616_t1, N3558);
nand NAND2_1123 (N3737, N3696, N3632);
nand NAND2_1124 (N3740, N3697, N3633);
nand NAND2_1125 (N3741, N3394_t1, N3716);
nand NAND2_1126 (N3742, N3397_t1, N3718);
nand NAND2_1127 (N3743, N3720, N3662);
and AND4_1128 (N3744, N3640_t0, N3647, N3644_t0, N3635_t0);
and AND2_1129 (N3745, N3635_t1, N3306);
and AND3_1130 (N3746, N3640_t1, N3635_t2, N3308);
and AND4_1131 (N3747, N3644_t1, N3635_t3, N3309, N3640_t2);
and AND2_1132 (N3748, N3648_t0, N3314);
and AND3_1133 (N3749, N3654_t0, N3648_t1, N3569);
not NOT1_1134 (N3750, N3721);
and AND2_1135 (N3753, N3722, N246_t5);
nand NAND2_1136 (N3754, N3728, N3692);
nand NAND2_1137 (N3758, N3729, N3694);
not NOT1_1138 (N3761, N3731);
or OR4_1139 (N3762, N3291, N3732, N3733, N3734);
nand NAND2_1140 (N3767, N3741, N3717);
nand NAND2_1141 (N3771, N3742, N3719);
not NOT1_1142 (N3774, N3744);
or OR4_1143 (N3775, N3304, N3745, N3746, N3747);
and AND2_1144 (N3778, N3723_t0, N3480);
and AND3_1145 (N3779, N3726, N3723_t1, N3409);
or OR2_1146 (N3780, N2125, N3753);
and AND2_1147 (N3790, N3750, N800_t1);
and AND2_1148 (N3793, N3737_t0, N3500);
and AND3_1149 (N3794, N3740, N3737_t1, N3428);
or OR3_1150 (N3802, N3479, N3778, N3779);
buf BUFF1_1151 (N3803, N3780_t0);
buf BUFF1_1152 (N3804, N3780_t1);
not NOT1_1153 (N3805, N3762_t0);
and AND5_1154 (N3806, N3622_t1, N3730, N3754_t0, N3616_t2, N3758_t0);
and AND4_1155 (N3807, N3754_t1, N3616_t3, N3559, N3622_t2);
and AND5_1156 (N3808, N3758_t1, N3754_t2, N3616_t4, N3498, N3622_t3);
buf BUFF1_1157 (N3809, N3790_t0);
or OR3_1158 (N3811, N3499, N3793, N3794);
not NOT1_1159 (N3812, N3775_t0);
and AND5_1160 (N3813, N3654_t1, N3743, N3767_t0, N3648_t2, N3771_t0);
and AND4_1161 (N3814, N3767_t1, N3648_t3, N3570, N3654_t2);
and AND5_1162 (N3815, N3771_t1, N3767_t2, N3648_t4, N3517, N3654_t3);
or OR5_1163 (N3816, N3299, N3735, N3736, N3807, N3808);
and AND2_1164 (N3817, N3806, N3802);
nand NAND2_1165 (N3818, N3805, N3761);
not NOT1_1166 (N3819, N3790_t1);
or OR5_1167 (N3820, N3312, N3748, N3749, N3814, N3815);
and AND2_1168 (N3821, N3813, N3811);
nand NAND2_1169 (N3822, N3812, N3774);
or OR2_1170 (N3823, N3816, N3817);
and AND3_1171 (N3826, N3727, N3819, N2841_t1);
or OR2_1172 (N3827, N3820, N3821);
not NOT1_1173 (N3834, N3823_t0);
and AND2_1174 (N3835, N3818, N3823_t1);
not NOT1_1175 (N3836, N3827_t0);
and AND2_1176 (N3837, N3822, N3827_t1);
and AND2_1177 (N3838, N3762_t1, N3834);
and AND2_1178 (N3839, N3775_t1, N3836);
or OR2_1179 (N3840, N3838, N3835);
or OR2_1180 (N3843, N3839, N3837);
buf BUFF1_1181 (N3851, N3843_t0);
nand NAND2_1182 (N3852, N3843_t1, N3840_t0);
and AND2_1183 (N3857, N3843_t2, N3852_t0);
and AND2_1184 (N3858, N3852_t1, N3840_t1);
or OR2_1185 (N3859, N3857, N3858);
not NOT1_1186 (N3864, N3859_t0);
and AND2_1187 (N3869, N3859_t1, N3864_t0);
or OR2_1188 (N3870, N3869, N3864_t1);
not NOT1_1189 (N3875, N3870_t0);
and AND3_1190 (N3876, N2826_t1, N3028, N3870_t1);
and AND3_1191 (N3877, N3826, N3876, N1591_t3);
buf BUFF1_1192 (N3881, N3877_t0);
not NOT1_1193 (N3882, N3877_t1);
buf BUFF1_1194 (N143_O, N143_I_t);
buf BUFF1_1195 (N144_O, N144_I_t);
buf BUFF1_1196 (N145_O, N145_I_t);
buf BUFF1_1197 (N146_O, N146_I_t);
buf BUFF1_1198 (N147_O, N147_I_t);
buf BUFF1_1199 (N148_O, N148_I_t);
buf BUFF1_1200 (N149_O, N149_I_t);
buf BUFF1_1201 (N150_O, N150_I_t);
buf BUFF1_1202 (N151_O, N151_I_t);
buf BUFF1_1203 (N152_O, N152_I_t);
buf BUFF1_1204 (N153_O, N153_I_t);
buf BUFF1_1205 (N154_O, N154_I_t);
buf BUFF1_1206 (N155_O, N155_I_t);
buf BUFF1_1207 (N156_O, N156_I_t);
buf BUFF1_1208 (N157_O, N157_I_t);
buf BUFF1_1209 (N158_O, N158_I_t);
buf BUFF1_1210 (N159_O, N159_I_t);
buf BUFF1_1211 (N160_O, N160_I_t);
buf BUFF1_1212 (N161_O, N161_I_t);
buf BUFF1_1213 (N162_O, N162_I_t);
buf BUFF1_1214 (N163_O, N163_I_t);
buf BUFF1_1215 (N164_O, N164_I_t);
buf BUFF1_1216 (N165_O, N165_I_t);
buf BUFF1_1217 (N166_O, N166_I_t);
buf BUFF1_1218 (N167_O, N167_I_t);
buf BUFF1_1219 (N168_O, N168_I_t);
buf BUFF1_1220 (N169_O, N169_I_t);
buf BUFF1_1221 (N170_O, N170_I_t);
buf BUFF1_1222 (N171_O, N171_I_t);
buf BUFF1_1223 (N172_O, N172_I_t);
buf BUFF1_1224 (N173_O, N173_I_t);
buf BUFF1_1225 (N174_O, N174_I_t);
buf BUFF1_1226 (N175_O, N175_I_t);
buf BUFF1_1227 (N176_O, N176_I_t);
buf BUFF1_1228 (N177_O, N177_I_t);
buf BUFF1_1229 (N178_O, N178_I_t);
buf BUFF1_1230 (N179_O, N179_I_t);
buf BUFF1_1231 (N180_O, N180_I_t);
buf BUFF1_1232 (N181_O, N181_I_t);
buf BUFF1_1233 (N182_O, N182_I_t);
buf BUFF1_1234 (N183_O, N183_I_t);
buf BUFF1_1235 (N184_O, N184_I_t);
buf BUFF1_1236 (N185_O, N185_I_t);
buf BUFF1_1237 (N186_O, N186_I_t);
buf BUFF1_1238 (N187_O, N187_I_t);
buf BUFF1_1239 (N188_O, N188_I_t);
buf BUFF1_1240 (N189_O, N189_I_t);
buf BUFF1_1241 (N190_O, N190_I_t);
buf BUFF1_1242 (N191_O, N191_I_t);
buf BUFF1_1243 (N192_O, N192_I_t);
buf BUFF1_1244 (N193_O, N193_I_t);
buf BUFF1_1245 (N194_O, N194_I_t);
buf BUFF1_1246 (N195_O, N195_I_t);
buf BUFF1_1247 (N196_O, N196_I_t);
buf BUFF1_1248 (N197_O, N197_I_t);
buf BUFF1_1249 (N198_O, N198_I_t);
buf BUFF1_1250 (N199_O, N199_I_t);
buf BUFF1_1251 (N200_O, N200_I_t);
buf BUFF1_1252 (N201_O, N201_I_t);
buf BUFF1_1253 (N202_O, N202_I_t);
buf BUFF1_1254 (N203_O, N203_I_t);
buf BUFF1_1255 (N204_O, N204_I_t);
buf BUFF1_1256 (N205_O, N205_I_t);
buf BUFF1_1257 (N206_O, N206_I_t);
buf BUFF1_1258 (N207_O, N207_I_t);
buf BUFF1_1259 (N208_O, N208_I_t);
buf BUFF1_1260 (N209_O, N209_I_t);
buf BUFF1_1261 (N210_O, N210_I_t);
buf BUFF1_1262 (N211_O, N211_I_t);
buf BUFF1_1263 (N212_O, N212_I_t);
buf BUFF1_1264 (N213_O, N213_I_t);
buf BUFF1_1265 (N214_O, N214_I_t);
buf BUFF1_1266 (N215_O, N215_I_t);
buf BUFF1_1267 (N216_O, N216_I_t);
buf BUFF1_1268 (N217_O, N217_I_t);
buf BUFF1_1269 (N218_O, N218_I_t);

endmodule
