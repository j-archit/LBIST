// ORA #1 - Result Compressor 

module rc
#(parameter OUTPUT_BITS = 4)
(
    input clk
);
    
endmodule