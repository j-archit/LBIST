/*
    Device Mid Section
    Consists of
        1. Fault Injection Logic (FIL)
        2. CUT - For Fault Injection
        3. CUT - Fault Free CUT

    Parameters:
        1. IN_BITS  : Number of Inputs / Input Bits
        2. OUT_BITS : Number of Outputs / Output Bits

    Inputs:
        1. clk      : Synchronizing Clock Input
        2. rst      : Asynch Reset (For FIL only)
        3. inc      : FIC Increment Signal (FIL injects New Fault in CUT when inc goes High)
        3. TEST_IP  : Input Test Pattern

    Outputs:
        1. CUT_OP   : Faulty Circuit Output
        2. FF_OP    : Fault Free Output

    Architecture:
        FIL, CUT1 and CUT2 are placed parallel, TEST_IP is given to both the CUTs. 
*/

`timescale 1ns/1ns

module mid
#(parameter IN_BITS = 1, parameter OUT_BITS = 1) 
(
    input clk,
    input rst,
    input FIL_INC,
    output FIL_END,
    input [IN_BITS-1:0] TEST_IP,
    output [OUT_BITS-1:0] CUT_OP, FF_OP
);
    
    // Python Script makes changes using "// Anchor" Comment
    // Make NO CHANGES in this block manually
    // Anchor
	c2670f #() faulty(
		FIL_INC, FIL_END, clk, rst, TEST_IP[232], TEST_IP[231], TEST_IP[230], TEST_IP[229], TEST_IP[228], TEST_IP[227], TEST_IP[226], TEST_IP[225], TEST_IP[224], TEST_IP[223], TEST_IP[222], TEST_IP[221], TEST_IP[220], TEST_IP[219], TEST_IP[218], TEST_IP[217], TEST_IP[216], TEST_IP[215], TEST_IP[214], TEST_IP[213], TEST_IP[212], TEST_IP[211], TEST_IP[210], TEST_IP[209], TEST_IP[208], TEST_IP[207], TEST_IP[206], TEST_IP[205], TEST_IP[204], TEST_IP[203], TEST_IP[202], TEST_IP[201], TEST_IP[200], TEST_IP[199], TEST_IP[198], TEST_IP[197], TEST_IP[196], TEST_IP[195], TEST_IP[194], TEST_IP[193], TEST_IP[192], TEST_IP[191], TEST_IP[190], TEST_IP[189], TEST_IP[188], TEST_IP[187], TEST_IP[186], TEST_IP[185], TEST_IP[184], TEST_IP[183], TEST_IP[182], TEST_IP[181], TEST_IP[180], TEST_IP[179], TEST_IP[178], TEST_IP[177], TEST_IP[176], TEST_IP[175], TEST_IP[174], TEST_IP[173], TEST_IP[172], TEST_IP[171], TEST_IP[170], TEST_IP[169], TEST_IP[168], TEST_IP[167], TEST_IP[166], TEST_IP[165], TEST_IP[164], TEST_IP[163], TEST_IP[162], TEST_IP[161], TEST_IP[160], TEST_IP[159], TEST_IP[158], TEST_IP[157], TEST_IP[156], TEST_IP[155], TEST_IP[154], TEST_IP[153], TEST_IP[152], TEST_IP[151], TEST_IP[150], TEST_IP[149], TEST_IP[148], TEST_IP[147], TEST_IP[146], TEST_IP[145], TEST_IP[144], TEST_IP[143], TEST_IP[142], TEST_IP[141], TEST_IP[140], TEST_IP[139], TEST_IP[138], TEST_IP[137], TEST_IP[136], TEST_IP[135], TEST_IP[134], TEST_IP[133], TEST_IP[132], TEST_IP[131], TEST_IP[130], TEST_IP[129], TEST_IP[128], TEST_IP[127], TEST_IP[126], TEST_IP[125], TEST_IP[124], TEST_IP[123], TEST_IP[122], TEST_IP[121], TEST_IP[120], TEST_IP[119], TEST_IP[118], TEST_IP[117], TEST_IP[116], TEST_IP[115], TEST_IP[114], TEST_IP[113], TEST_IP[112], TEST_IP[111], TEST_IP[110], TEST_IP[109], TEST_IP[108], TEST_IP[107], TEST_IP[106], TEST_IP[105], TEST_IP[104], TEST_IP[103], TEST_IP[102], TEST_IP[101], TEST_IP[100], TEST_IP[99], TEST_IP[98], TEST_IP[97], TEST_IP[96], TEST_IP[95], TEST_IP[94], TEST_IP[93], TEST_IP[92], TEST_IP[91], TEST_IP[90], TEST_IP[89], TEST_IP[88], TEST_IP[87], TEST_IP[86], TEST_IP[85], TEST_IP[84], TEST_IP[83], TEST_IP[82], TEST_IP[81], TEST_IP[80], TEST_IP[79], TEST_IP[78], TEST_IP[77], TEST_IP[76], TEST_IP[75], TEST_IP[74], TEST_IP[73], TEST_IP[72], TEST_IP[71], TEST_IP[70], TEST_IP[69], TEST_IP[68], TEST_IP[67], TEST_IP[66], TEST_IP[65], TEST_IP[64], TEST_IP[63], TEST_IP[62], TEST_IP[61], TEST_IP[60], TEST_IP[59], TEST_IP[58], TEST_IP[57], TEST_IP[56], TEST_IP[55], TEST_IP[54], TEST_IP[53], TEST_IP[52], TEST_IP[51], TEST_IP[50], TEST_IP[49], TEST_IP[48], TEST_IP[47], TEST_IP[46], TEST_IP[45], TEST_IP[44], TEST_IP[43], TEST_IP[42], TEST_IP[41], TEST_IP[40], TEST_IP[39], TEST_IP[38], TEST_IP[37], TEST_IP[36], TEST_IP[35], TEST_IP[34], TEST_IP[33], TEST_IP[32], TEST_IP[31], TEST_IP[30], TEST_IP[29], TEST_IP[28], TEST_IP[27], TEST_IP[26], TEST_IP[25], TEST_IP[24], TEST_IP[23], TEST_IP[22], TEST_IP[21], TEST_IP[20], TEST_IP[19], TEST_IP[18], TEST_IP[17], TEST_IP[16], TEST_IP[15], TEST_IP[14], TEST_IP[13], TEST_IP[12], TEST_IP[11], TEST_IP[10], TEST_IP[9], TEST_IP[8], TEST_IP[7], TEST_IP[6], TEST_IP[5], TEST_IP[4], TEST_IP[3], TEST_IP[2], TEST_IP[1], TEST_IP[0], CUT_OP[139], CUT_OP[138], CUT_OP[137], CUT_OP[136], CUT_OP[135], CUT_OP[134], CUT_OP[133], CUT_OP[132], CUT_OP[131], CUT_OP[130], CUT_OP[129], CUT_OP[128], CUT_OP[127], CUT_OP[126], CUT_OP[125], CUT_OP[124], CUT_OP[123], CUT_OP[122], CUT_OP[121], CUT_OP[120], CUT_OP[119], CUT_OP[118], CUT_OP[117], CUT_OP[116], CUT_OP[115], CUT_OP[114], CUT_OP[113], CUT_OP[112], CUT_OP[111], CUT_OP[110], CUT_OP[109], CUT_OP[108], CUT_OP[107], CUT_OP[106], CUT_OP[105], CUT_OP[104], CUT_OP[103], CUT_OP[102], CUT_OP[101], CUT_OP[100], CUT_OP[99], CUT_OP[98], CUT_OP[97], CUT_OP[96], CUT_OP[95], CUT_OP[94], CUT_OP[93], CUT_OP[92], CUT_OP[91], CUT_OP[90], CUT_OP[89], CUT_OP[88], CUT_OP[87], CUT_OP[86], CUT_OP[85], CUT_OP[84], CUT_OP[83], CUT_OP[82], CUT_OP[81], CUT_OP[80], CUT_OP[79], CUT_OP[78], CUT_OP[77], CUT_OP[76], CUT_OP[75], CUT_OP[74], CUT_OP[73], CUT_OP[72], CUT_OP[71], CUT_OP[70], CUT_OP[69], CUT_OP[68], CUT_OP[67], CUT_OP[66], CUT_OP[65], CUT_OP[64], CUT_OP[63], CUT_OP[62], CUT_OP[61], CUT_OP[60], CUT_OP[59], CUT_OP[58], CUT_OP[57], CUT_OP[56], CUT_OP[55], CUT_OP[54], CUT_OP[53], CUT_OP[52], CUT_OP[51], CUT_OP[50], CUT_OP[49], CUT_OP[48], CUT_OP[47], CUT_OP[46], CUT_OP[45], CUT_OP[44], CUT_OP[43], CUT_OP[42], CUT_OP[41], CUT_OP[40], CUT_OP[39], CUT_OP[38], CUT_OP[37], CUT_OP[36], CUT_OP[35], CUT_OP[34], CUT_OP[33], CUT_OP[32], CUT_OP[31], CUT_OP[30], CUT_OP[29], CUT_OP[28], CUT_OP[27], CUT_OP[26], CUT_OP[25], CUT_OP[24], CUT_OP[23], CUT_OP[22], CUT_OP[21], CUT_OP[20], CUT_OP[19], CUT_OP[18], CUT_OP[17], CUT_OP[16], CUT_OP[15], CUT_OP[14], CUT_OP[13], CUT_OP[12], CUT_OP[11], CUT_OP[10], CUT_OP[9], CUT_OP[8], CUT_OP[7], CUT_OP[6], CUT_OP[5], CUT_OP[4], CUT_OP[3], CUT_OP[2], CUT_OP[1], CUT_OP[0]
    );
	c2670 #() faultf(
		TEST_IP[232], TEST_IP[231], TEST_IP[230], TEST_IP[229], TEST_IP[228], TEST_IP[227], TEST_IP[226], TEST_IP[225], TEST_IP[224], TEST_IP[223], TEST_IP[222], TEST_IP[221], TEST_IP[220], TEST_IP[219], TEST_IP[218], TEST_IP[217], TEST_IP[216], TEST_IP[215], TEST_IP[214], TEST_IP[213], TEST_IP[212], TEST_IP[211], TEST_IP[210], TEST_IP[209], TEST_IP[208], TEST_IP[207], TEST_IP[206], TEST_IP[205], TEST_IP[204], TEST_IP[203], TEST_IP[202], TEST_IP[201], TEST_IP[200], TEST_IP[199], TEST_IP[198], TEST_IP[197], TEST_IP[196], TEST_IP[195], TEST_IP[194], TEST_IP[193], TEST_IP[192], TEST_IP[191], TEST_IP[190], TEST_IP[189], TEST_IP[188], TEST_IP[187], TEST_IP[186], TEST_IP[185], TEST_IP[184], TEST_IP[183], TEST_IP[182], TEST_IP[181], TEST_IP[180], TEST_IP[179], TEST_IP[178], TEST_IP[177], TEST_IP[176], TEST_IP[175], TEST_IP[174], TEST_IP[173], TEST_IP[172], TEST_IP[171], TEST_IP[170], TEST_IP[169], TEST_IP[168], TEST_IP[167], TEST_IP[166], TEST_IP[165], TEST_IP[164], TEST_IP[163], TEST_IP[162], TEST_IP[161], TEST_IP[160], TEST_IP[159], TEST_IP[158], TEST_IP[157], TEST_IP[156], TEST_IP[155], TEST_IP[154], TEST_IP[153], TEST_IP[152], TEST_IP[151], TEST_IP[150], TEST_IP[149], TEST_IP[148], TEST_IP[147], TEST_IP[146], TEST_IP[145], TEST_IP[144], TEST_IP[143], TEST_IP[142], TEST_IP[141], TEST_IP[140], TEST_IP[139], TEST_IP[138], TEST_IP[137], TEST_IP[136], TEST_IP[135], TEST_IP[134], TEST_IP[133], TEST_IP[132], TEST_IP[131], TEST_IP[130], TEST_IP[129], TEST_IP[128], TEST_IP[127], TEST_IP[126], TEST_IP[125], TEST_IP[124], TEST_IP[123], TEST_IP[122], TEST_IP[121], TEST_IP[120], TEST_IP[119], TEST_IP[118], TEST_IP[117], TEST_IP[116], TEST_IP[115], TEST_IP[114], TEST_IP[113], TEST_IP[112], TEST_IP[111], TEST_IP[110], TEST_IP[109], TEST_IP[108], TEST_IP[107], TEST_IP[106], TEST_IP[105], TEST_IP[104], TEST_IP[103], TEST_IP[102], TEST_IP[101], TEST_IP[100], TEST_IP[99], TEST_IP[98], TEST_IP[97], TEST_IP[96], TEST_IP[95], TEST_IP[94], TEST_IP[93], TEST_IP[92], TEST_IP[91], TEST_IP[90], TEST_IP[89], TEST_IP[88], TEST_IP[87], TEST_IP[86], TEST_IP[85], TEST_IP[84], TEST_IP[83], TEST_IP[82], TEST_IP[81], TEST_IP[80], TEST_IP[79], TEST_IP[78], TEST_IP[77], TEST_IP[76], TEST_IP[75], TEST_IP[74], TEST_IP[73], TEST_IP[72], TEST_IP[71], TEST_IP[70], TEST_IP[69], TEST_IP[68], TEST_IP[67], TEST_IP[66], TEST_IP[65], TEST_IP[64], TEST_IP[63], TEST_IP[62], TEST_IP[61], TEST_IP[60], TEST_IP[59], TEST_IP[58], TEST_IP[57], TEST_IP[56], TEST_IP[55], TEST_IP[54], TEST_IP[53], TEST_IP[52], TEST_IP[51], TEST_IP[50], TEST_IP[49], TEST_IP[48], TEST_IP[47], TEST_IP[46], TEST_IP[45], TEST_IP[44], TEST_IP[43], TEST_IP[42], TEST_IP[41], TEST_IP[40], TEST_IP[39], TEST_IP[38], TEST_IP[37], TEST_IP[36], TEST_IP[35], TEST_IP[34], TEST_IP[33], TEST_IP[32], TEST_IP[31], TEST_IP[30], TEST_IP[29], TEST_IP[28], TEST_IP[27], TEST_IP[26], TEST_IP[25], TEST_IP[24], TEST_IP[23], TEST_IP[22], TEST_IP[21], TEST_IP[20], TEST_IP[19], TEST_IP[18], TEST_IP[17], TEST_IP[16], TEST_IP[15], TEST_IP[14], TEST_IP[13], TEST_IP[12], TEST_IP[11], TEST_IP[10], TEST_IP[9], TEST_IP[8], TEST_IP[7], TEST_IP[6], TEST_IP[5], TEST_IP[4], TEST_IP[3], TEST_IP[2], TEST_IP[1], TEST_IP[0], FF_OP[139], FF_OP[138], FF_OP[137], FF_OP[136], FF_OP[135], FF_OP[134], FF_OP[133], FF_OP[132], FF_OP[131], FF_OP[130], FF_OP[129], FF_OP[128], FF_OP[127], FF_OP[126], FF_OP[125], FF_OP[124], FF_OP[123], FF_OP[122], FF_OP[121], FF_OP[120], FF_OP[119], FF_OP[118], FF_OP[117], FF_OP[116], FF_OP[115], FF_OP[114], FF_OP[113], FF_OP[112], FF_OP[111], FF_OP[110], FF_OP[109], FF_OP[108], FF_OP[107], FF_OP[106], FF_OP[105], FF_OP[104], FF_OP[103], FF_OP[102], FF_OP[101], FF_OP[100], FF_OP[99], FF_OP[98], FF_OP[97], FF_OP[96], FF_OP[95], FF_OP[94], FF_OP[93], FF_OP[92], FF_OP[91], FF_OP[90], FF_OP[89], FF_OP[88], FF_OP[87], FF_OP[86], FF_OP[85], FF_OP[84], FF_OP[83], FF_OP[82], FF_OP[81], FF_OP[80], FF_OP[79], FF_OP[78], FF_OP[77], FF_OP[76], FF_OP[75], FF_OP[74], FF_OP[73], FF_OP[72], FF_OP[71], FF_OP[70], FF_OP[69], FF_OP[68], FF_OP[67], FF_OP[66], FF_OP[65], FF_OP[64], FF_OP[63], FF_OP[62], FF_OP[61], FF_OP[60], FF_OP[59], FF_OP[58], FF_OP[57], FF_OP[56], FF_OP[55], FF_OP[54], FF_OP[53], FF_OP[52], FF_OP[51], FF_OP[50], FF_OP[49], FF_OP[48], FF_OP[47], FF_OP[46], FF_OP[45], FF_OP[44], FF_OP[43], FF_OP[42], FF_OP[41], FF_OP[40], FF_OP[39], FF_OP[38], FF_OP[37], FF_OP[36], FF_OP[35], FF_OP[34], FF_OP[33], FF_OP[32], FF_OP[31], FF_OP[30], FF_OP[29], FF_OP[28], FF_OP[27], FF_OP[26], FF_OP[25], FF_OP[24], FF_OP[23], FF_OP[22], FF_OP[21], FF_OP[20], FF_OP[19], FF_OP[18], FF_OP[17], FF_OP[16], FF_OP[15], FF_OP[14], FF_OP[13], FF_OP[12], FF_OP[11], FF_OP[10], FF_OP[9], FF_OP[8], FF_OP[7], FF_OP[6], FF_OP[5], FF_OP[4], FF_OP[3], FF_OP[2], FF_OP[1], FF_OP[0]
    );
    // Block Ends
    
endmodule