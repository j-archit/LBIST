// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8
// Nfaults 528

`timescale 1ns/1ns

module c499f (INC,END,clk,rst,N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

// FaultModel
input INC,clk,rst;
output reg END;
reg fault;
wire N129_t,N130_t,N131_t,N132_t,N133_t,N134_t,N135_t,N136_t;
wire N1_t0,N1_t1,N1_t2,N5_t0,N5_t1,N5_t2,N9_t0,N9_t1,N9_t2,
     N13_t0,N13_t1,N13_t2,N17_t0,N17_t1,N17_t2,N21_t0,N21_t1,N21_t2,N25_t0,
     N25_t1,N25_t2,N29_t0,N29_t1,N29_t2,N33_t0,N33_t1,N33_t2,N37_t0,N37_t1,
     N37_t2,N41_t0,N41_t1,N41_t2,N45_t0,N45_t1,N45_t2,N49_t0,N49_t1,N49_t2,
     N53_t0,N53_t1,N53_t2,N57_t0,N57_t1,N57_t2,N61_t0,N61_t1,N61_t2,N65_t0,
     N65_t1,N65_t2,N69_t0,N69_t1,N69_t2,N73_t0,N73_t1,N73_t2,N77_t0,N77_t1,
     N77_t2,N81_t0,N81_t1,N81_t2,N85_t0,N85_t1,N85_t2,N89_t0,N89_t1,N89_t2,
     N93_t0,N93_t1,N93_t2,N97_t0,N97_t1,N97_t2,N101_t0,N101_t1,N101_t2,N105_t0,
     N105_t1,N105_t2,N109_t0,N109_t1,N109_t2,N113_t0,N113_t1,N113_t2,N117_t0,N117_t1,
     N117_t2,N121_t0,N121_t1,N121_t2,N125_t0,N125_t1,N125_t2,N137_t0,N137_t1,N137_t2,
     N137_t3,N137_t4,N137_t5,N137_t6,N137_t7,N290_t0,N290_t1,N293_t0,N293_t1,N296_t0,
     N296_t1,N299_t0,N299_t1,N302_t0,N302_t1,N305_t0,N305_t1,N308_t0,N308_t1,N311_t0,
     N311_t1,N354_t0,N354_t1,N354_t2,N354_t3,N354_t4,N354_t5,N354_t6,N354_t7,N354_t8,
     N354_t9,N354_t10,N354_t11,N367_t0,N367_t1,N367_t2,N367_t3,N367_t4,N367_t5,N367_t6,
     N367_t7,N367_t8,N367_t9,N367_t10,N367_t11,N380_t0,N380_t1,N380_t2,N380_t3,N380_t4,
     N380_t5,N380_t6,N380_t7,N380_t8,N380_t9,N380_t10,N380_t11,N393_t0,N393_t1,N393_t2,
     N393_t3,N393_t4,N393_t5,N393_t6,N393_t7,N393_t8,N393_t9,N393_t10,N393_t11,N419_t0,
     N419_t1,N419_t2,N419_t3,N419_t4,N419_t5,N419_t6,N419_t7,N419_t8,N419_t9,N419_t10,
     N419_t11,N445_t0,N445_t1,N445_t2,N445_t3,N445_t4,N445_t5,N445_t6,N445_t7,N445_t8,
     N445_t9,N445_t10,N445_t11,N432_t0,N432_t1,N432_t2,N432_t3,N432_t4,N432_t5,N432_t6,
     N432_t7,N432_t8,N432_t9,N432_t10,N432_t11,N406_t0,N406_t1,N406_t2,N406_t3,N406_t4,
     N406_t5,N406_t6,N406_t7,N406_t8,N406_t9,N406_t10,N406_t11,N602_t0,N602_t1,N602_t2,
     N602_t3,N607_t0,N607_t1,N607_t2,N607_t3,N620_t0,N620_t1,N620_t2,N620_t3,N625_t0,
     N625_t1,N625_t2,N625_t3,N630_t0,N630_t1,N630_t2,N630_t3,N635_t0,N635_t1,N635_t2,
     N635_t3,N640_t0,N640_t1,N640_t2,N640_t3,N645_t0,N645_t1,N645_t2,N645_t3,N650_t0,
     N650_t1,N650_t2,N650_t3,N655_t0,N655_t1,N655_t2,N655_t3;
reg [263:0] FEN;
fim PI_N129( .fault(fault), .net(N129), .FEN(FEN[0]), .op(N129_t) );
fim PI_N130( .fault(fault), .net(N130), .FEN(FEN[1]), .op(N130_t) );
fim PI_N131( .fault(fault), .net(N131), .FEN(FEN[2]), .op(N131_t) );
fim PI_N132( .fault(fault), .net(N132), .FEN(FEN[3]), .op(N132_t) );
fim PI_N133( .fault(fault), .net(N133), .FEN(FEN[4]), .op(N133_t) );
fim PI_N134( .fault(fault), .net(N134), .FEN(FEN[5]), .op(N134_t) );
fim PI_N135( .fault(fault), .net(N135), .FEN(FEN[6]), .op(N135_t) );
fim PI_N136( .fault(fault), .net(N136), .FEN(FEN[7]), .op(N136_t) );
fim FAN_N1_0 ( .fault(fault), .net(N1), .FEN(FEN[8]), .op(N1_t0) );
fim FAN_N1_1 ( .fault(fault), .net(N1), .FEN(FEN[9]), .op(N1_t1) );
fim FAN_N1_2 ( .fault(fault), .net(N1), .FEN(FEN[10]), .op(N1_t2) );
fim FAN_N5_0 ( .fault(fault), .net(N5), .FEN(FEN[11]), .op(N5_t0) );
fim FAN_N5_1 ( .fault(fault), .net(N5), .FEN(FEN[12]), .op(N5_t1) );
fim FAN_N5_2 ( .fault(fault), .net(N5), .FEN(FEN[13]), .op(N5_t2) );
fim FAN_N9_0 ( .fault(fault), .net(N9), .FEN(FEN[14]), .op(N9_t0) );
fim FAN_N9_1 ( .fault(fault), .net(N9), .FEN(FEN[15]), .op(N9_t1) );
fim FAN_N9_2 ( .fault(fault), .net(N9), .FEN(FEN[16]), .op(N9_t2) );
fim FAN_N13_0 ( .fault(fault), .net(N13), .FEN(FEN[17]), .op(N13_t0) );
fim FAN_N13_1 ( .fault(fault), .net(N13), .FEN(FEN[18]), .op(N13_t1) );
fim FAN_N13_2 ( .fault(fault), .net(N13), .FEN(FEN[19]), .op(N13_t2) );
fim FAN_N17_0 ( .fault(fault), .net(N17), .FEN(FEN[20]), .op(N17_t0) );
fim FAN_N17_1 ( .fault(fault), .net(N17), .FEN(FEN[21]), .op(N17_t1) );
fim FAN_N17_2 ( .fault(fault), .net(N17), .FEN(FEN[22]), .op(N17_t2) );
fim FAN_N21_0 ( .fault(fault), .net(N21), .FEN(FEN[23]), .op(N21_t0) );
fim FAN_N21_1 ( .fault(fault), .net(N21), .FEN(FEN[24]), .op(N21_t1) );
fim FAN_N21_2 ( .fault(fault), .net(N21), .FEN(FEN[25]), .op(N21_t2) );
fim FAN_N25_0 ( .fault(fault), .net(N25), .FEN(FEN[26]), .op(N25_t0) );
fim FAN_N25_1 ( .fault(fault), .net(N25), .FEN(FEN[27]), .op(N25_t1) );
fim FAN_N25_2 ( .fault(fault), .net(N25), .FEN(FEN[28]), .op(N25_t2) );
fim FAN_N29_0 ( .fault(fault), .net(N29), .FEN(FEN[29]), .op(N29_t0) );
fim FAN_N29_1 ( .fault(fault), .net(N29), .FEN(FEN[30]), .op(N29_t1) );
fim FAN_N29_2 ( .fault(fault), .net(N29), .FEN(FEN[31]), .op(N29_t2) );
fim FAN_N33_0 ( .fault(fault), .net(N33), .FEN(FEN[32]), .op(N33_t0) );
fim FAN_N33_1 ( .fault(fault), .net(N33), .FEN(FEN[33]), .op(N33_t1) );
fim FAN_N33_2 ( .fault(fault), .net(N33), .FEN(FEN[34]), .op(N33_t2) );
fim FAN_N37_0 ( .fault(fault), .net(N37), .FEN(FEN[35]), .op(N37_t0) );
fim FAN_N37_1 ( .fault(fault), .net(N37), .FEN(FEN[36]), .op(N37_t1) );
fim FAN_N37_2 ( .fault(fault), .net(N37), .FEN(FEN[37]), .op(N37_t2) );
fim FAN_N41_0 ( .fault(fault), .net(N41), .FEN(FEN[38]), .op(N41_t0) );
fim FAN_N41_1 ( .fault(fault), .net(N41), .FEN(FEN[39]), .op(N41_t1) );
fim FAN_N41_2 ( .fault(fault), .net(N41), .FEN(FEN[40]), .op(N41_t2) );
fim FAN_N45_0 ( .fault(fault), .net(N45), .FEN(FEN[41]), .op(N45_t0) );
fim FAN_N45_1 ( .fault(fault), .net(N45), .FEN(FEN[42]), .op(N45_t1) );
fim FAN_N45_2 ( .fault(fault), .net(N45), .FEN(FEN[43]), .op(N45_t2) );
fim FAN_N49_0 ( .fault(fault), .net(N49), .FEN(FEN[44]), .op(N49_t0) );
fim FAN_N49_1 ( .fault(fault), .net(N49), .FEN(FEN[45]), .op(N49_t1) );
fim FAN_N49_2 ( .fault(fault), .net(N49), .FEN(FEN[46]), .op(N49_t2) );
fim FAN_N53_0 ( .fault(fault), .net(N53), .FEN(FEN[47]), .op(N53_t0) );
fim FAN_N53_1 ( .fault(fault), .net(N53), .FEN(FEN[48]), .op(N53_t1) );
fim FAN_N53_2 ( .fault(fault), .net(N53), .FEN(FEN[49]), .op(N53_t2) );
fim FAN_N57_0 ( .fault(fault), .net(N57), .FEN(FEN[50]), .op(N57_t0) );
fim FAN_N57_1 ( .fault(fault), .net(N57), .FEN(FEN[51]), .op(N57_t1) );
fim FAN_N57_2 ( .fault(fault), .net(N57), .FEN(FEN[52]), .op(N57_t2) );
fim FAN_N61_0 ( .fault(fault), .net(N61), .FEN(FEN[53]), .op(N61_t0) );
fim FAN_N61_1 ( .fault(fault), .net(N61), .FEN(FEN[54]), .op(N61_t1) );
fim FAN_N61_2 ( .fault(fault), .net(N61), .FEN(FEN[55]), .op(N61_t2) );
fim FAN_N65_0 ( .fault(fault), .net(N65), .FEN(FEN[56]), .op(N65_t0) );
fim FAN_N65_1 ( .fault(fault), .net(N65), .FEN(FEN[57]), .op(N65_t1) );
fim FAN_N65_2 ( .fault(fault), .net(N65), .FEN(FEN[58]), .op(N65_t2) );
fim FAN_N69_0 ( .fault(fault), .net(N69), .FEN(FEN[59]), .op(N69_t0) );
fim FAN_N69_1 ( .fault(fault), .net(N69), .FEN(FEN[60]), .op(N69_t1) );
fim FAN_N69_2 ( .fault(fault), .net(N69), .FEN(FEN[61]), .op(N69_t2) );
fim FAN_N73_0 ( .fault(fault), .net(N73), .FEN(FEN[62]), .op(N73_t0) );
fim FAN_N73_1 ( .fault(fault), .net(N73), .FEN(FEN[63]), .op(N73_t1) );
fim FAN_N73_2 ( .fault(fault), .net(N73), .FEN(FEN[64]), .op(N73_t2) );
fim FAN_N77_0 ( .fault(fault), .net(N77), .FEN(FEN[65]), .op(N77_t0) );
fim FAN_N77_1 ( .fault(fault), .net(N77), .FEN(FEN[66]), .op(N77_t1) );
fim FAN_N77_2 ( .fault(fault), .net(N77), .FEN(FEN[67]), .op(N77_t2) );
fim FAN_N81_0 ( .fault(fault), .net(N81), .FEN(FEN[68]), .op(N81_t0) );
fim FAN_N81_1 ( .fault(fault), .net(N81), .FEN(FEN[69]), .op(N81_t1) );
fim FAN_N81_2 ( .fault(fault), .net(N81), .FEN(FEN[70]), .op(N81_t2) );
fim FAN_N85_0 ( .fault(fault), .net(N85), .FEN(FEN[71]), .op(N85_t0) );
fim FAN_N85_1 ( .fault(fault), .net(N85), .FEN(FEN[72]), .op(N85_t1) );
fim FAN_N85_2 ( .fault(fault), .net(N85), .FEN(FEN[73]), .op(N85_t2) );
fim FAN_N89_0 ( .fault(fault), .net(N89), .FEN(FEN[74]), .op(N89_t0) );
fim FAN_N89_1 ( .fault(fault), .net(N89), .FEN(FEN[75]), .op(N89_t1) );
fim FAN_N89_2 ( .fault(fault), .net(N89), .FEN(FEN[76]), .op(N89_t2) );
fim FAN_N93_0 ( .fault(fault), .net(N93), .FEN(FEN[77]), .op(N93_t0) );
fim FAN_N93_1 ( .fault(fault), .net(N93), .FEN(FEN[78]), .op(N93_t1) );
fim FAN_N93_2 ( .fault(fault), .net(N93), .FEN(FEN[79]), .op(N93_t2) );
fim FAN_N97_0 ( .fault(fault), .net(N97), .FEN(FEN[80]), .op(N97_t0) );
fim FAN_N97_1 ( .fault(fault), .net(N97), .FEN(FEN[81]), .op(N97_t1) );
fim FAN_N97_2 ( .fault(fault), .net(N97), .FEN(FEN[82]), .op(N97_t2) );
fim FAN_N101_0 ( .fault(fault), .net(N101), .FEN(FEN[83]), .op(N101_t0) );
fim FAN_N101_1 ( .fault(fault), .net(N101), .FEN(FEN[84]), .op(N101_t1) );
fim FAN_N101_2 ( .fault(fault), .net(N101), .FEN(FEN[85]), .op(N101_t2) );
fim FAN_N105_0 ( .fault(fault), .net(N105), .FEN(FEN[86]), .op(N105_t0) );
fim FAN_N105_1 ( .fault(fault), .net(N105), .FEN(FEN[87]), .op(N105_t1) );
fim FAN_N105_2 ( .fault(fault), .net(N105), .FEN(FEN[88]), .op(N105_t2) );
fim FAN_N109_0 ( .fault(fault), .net(N109), .FEN(FEN[89]), .op(N109_t0) );
fim FAN_N109_1 ( .fault(fault), .net(N109), .FEN(FEN[90]), .op(N109_t1) );
fim FAN_N109_2 ( .fault(fault), .net(N109), .FEN(FEN[91]), .op(N109_t2) );
fim FAN_N113_0 ( .fault(fault), .net(N113), .FEN(FEN[92]), .op(N113_t0) );
fim FAN_N113_1 ( .fault(fault), .net(N113), .FEN(FEN[93]), .op(N113_t1) );
fim FAN_N113_2 ( .fault(fault), .net(N113), .FEN(FEN[94]), .op(N113_t2) );
fim FAN_N117_0 ( .fault(fault), .net(N117), .FEN(FEN[95]), .op(N117_t0) );
fim FAN_N117_1 ( .fault(fault), .net(N117), .FEN(FEN[96]), .op(N117_t1) );
fim FAN_N117_2 ( .fault(fault), .net(N117), .FEN(FEN[97]), .op(N117_t2) );
fim FAN_N121_0 ( .fault(fault), .net(N121), .FEN(FEN[98]), .op(N121_t0) );
fim FAN_N121_1 ( .fault(fault), .net(N121), .FEN(FEN[99]), .op(N121_t1) );
fim FAN_N121_2 ( .fault(fault), .net(N121), .FEN(FEN[100]), .op(N121_t2) );
fim FAN_N125_0 ( .fault(fault), .net(N125), .FEN(FEN[101]), .op(N125_t0) );
fim FAN_N125_1 ( .fault(fault), .net(N125), .FEN(FEN[102]), .op(N125_t1) );
fim FAN_N125_2 ( .fault(fault), .net(N125), .FEN(FEN[103]), .op(N125_t2) );
fim FAN_N137_0 ( .fault(fault), .net(N137), .FEN(FEN[104]), .op(N137_t0) );
fim FAN_N137_1 ( .fault(fault), .net(N137), .FEN(FEN[105]), .op(N137_t1) );
fim FAN_N137_2 ( .fault(fault), .net(N137), .FEN(FEN[106]), .op(N137_t2) );
fim FAN_N137_3 ( .fault(fault), .net(N137), .FEN(FEN[107]), .op(N137_t3) );
fim FAN_N137_4 ( .fault(fault), .net(N137), .FEN(FEN[108]), .op(N137_t4) );
fim FAN_N137_5 ( .fault(fault), .net(N137), .FEN(FEN[109]), .op(N137_t5) );
fim FAN_N137_6 ( .fault(fault), .net(N137), .FEN(FEN[110]), .op(N137_t6) );
fim FAN_N137_7 ( .fault(fault), .net(N137), .FEN(FEN[111]), .op(N137_t7) );
fim FAN_N290_0 ( .fault(fault), .net(N290), .FEN(FEN[112]), .op(N290_t0) );
fim FAN_N290_1 ( .fault(fault), .net(N290), .FEN(FEN[113]), .op(N290_t1) );
fim FAN_N293_0 ( .fault(fault), .net(N293), .FEN(FEN[114]), .op(N293_t0) );
fim FAN_N293_1 ( .fault(fault), .net(N293), .FEN(FEN[115]), .op(N293_t1) );
fim FAN_N296_0 ( .fault(fault), .net(N296), .FEN(FEN[116]), .op(N296_t0) );
fim FAN_N296_1 ( .fault(fault), .net(N296), .FEN(FEN[117]), .op(N296_t1) );
fim FAN_N299_0 ( .fault(fault), .net(N299), .FEN(FEN[118]), .op(N299_t0) );
fim FAN_N299_1 ( .fault(fault), .net(N299), .FEN(FEN[119]), .op(N299_t1) );
fim FAN_N302_0 ( .fault(fault), .net(N302), .FEN(FEN[120]), .op(N302_t0) );
fim FAN_N302_1 ( .fault(fault), .net(N302), .FEN(FEN[121]), .op(N302_t1) );
fim FAN_N305_0 ( .fault(fault), .net(N305), .FEN(FEN[122]), .op(N305_t0) );
fim FAN_N305_1 ( .fault(fault), .net(N305), .FEN(FEN[123]), .op(N305_t1) );
fim FAN_N308_0 ( .fault(fault), .net(N308), .FEN(FEN[124]), .op(N308_t0) );
fim FAN_N308_1 ( .fault(fault), .net(N308), .FEN(FEN[125]), .op(N308_t1) );
fim FAN_N311_0 ( .fault(fault), .net(N311), .FEN(FEN[126]), .op(N311_t0) );
fim FAN_N311_1 ( .fault(fault), .net(N311), .FEN(FEN[127]), .op(N311_t1) );
fim FAN_N354_0 ( .fault(fault), .net(N354), .FEN(FEN[128]), .op(N354_t0) );
fim FAN_N354_1 ( .fault(fault), .net(N354), .FEN(FEN[129]), .op(N354_t1) );
fim FAN_N354_2 ( .fault(fault), .net(N354), .FEN(FEN[130]), .op(N354_t2) );
fim FAN_N354_3 ( .fault(fault), .net(N354), .FEN(FEN[131]), .op(N354_t3) );
fim FAN_N354_4 ( .fault(fault), .net(N354), .FEN(FEN[132]), .op(N354_t4) );
fim FAN_N354_5 ( .fault(fault), .net(N354), .FEN(FEN[133]), .op(N354_t5) );
fim FAN_N354_6 ( .fault(fault), .net(N354), .FEN(FEN[134]), .op(N354_t6) );
fim FAN_N354_7 ( .fault(fault), .net(N354), .FEN(FEN[135]), .op(N354_t7) );
fim FAN_N354_8 ( .fault(fault), .net(N354), .FEN(FEN[136]), .op(N354_t8) );
fim FAN_N354_9 ( .fault(fault), .net(N354), .FEN(FEN[137]), .op(N354_t9) );
fim FAN_N354_10 ( .fault(fault), .net(N354), .FEN(FEN[138]), .op(N354_t10) );
fim FAN_N354_11 ( .fault(fault), .net(N354), .FEN(FEN[139]), .op(N354_t11) );
fim FAN_N367_0 ( .fault(fault), .net(N367), .FEN(FEN[140]), .op(N367_t0) );
fim FAN_N367_1 ( .fault(fault), .net(N367), .FEN(FEN[141]), .op(N367_t1) );
fim FAN_N367_2 ( .fault(fault), .net(N367), .FEN(FEN[142]), .op(N367_t2) );
fim FAN_N367_3 ( .fault(fault), .net(N367), .FEN(FEN[143]), .op(N367_t3) );
fim FAN_N367_4 ( .fault(fault), .net(N367), .FEN(FEN[144]), .op(N367_t4) );
fim FAN_N367_5 ( .fault(fault), .net(N367), .FEN(FEN[145]), .op(N367_t5) );
fim FAN_N367_6 ( .fault(fault), .net(N367), .FEN(FEN[146]), .op(N367_t6) );
fim FAN_N367_7 ( .fault(fault), .net(N367), .FEN(FEN[147]), .op(N367_t7) );
fim FAN_N367_8 ( .fault(fault), .net(N367), .FEN(FEN[148]), .op(N367_t8) );
fim FAN_N367_9 ( .fault(fault), .net(N367), .FEN(FEN[149]), .op(N367_t9) );
fim FAN_N367_10 ( .fault(fault), .net(N367), .FEN(FEN[150]), .op(N367_t10) );
fim FAN_N367_11 ( .fault(fault), .net(N367), .FEN(FEN[151]), .op(N367_t11) );
fim FAN_N380_0 ( .fault(fault), .net(N380), .FEN(FEN[152]), .op(N380_t0) );
fim FAN_N380_1 ( .fault(fault), .net(N380), .FEN(FEN[153]), .op(N380_t1) );
fim FAN_N380_2 ( .fault(fault), .net(N380), .FEN(FEN[154]), .op(N380_t2) );
fim FAN_N380_3 ( .fault(fault), .net(N380), .FEN(FEN[155]), .op(N380_t3) );
fim FAN_N380_4 ( .fault(fault), .net(N380), .FEN(FEN[156]), .op(N380_t4) );
fim FAN_N380_5 ( .fault(fault), .net(N380), .FEN(FEN[157]), .op(N380_t5) );
fim FAN_N380_6 ( .fault(fault), .net(N380), .FEN(FEN[158]), .op(N380_t6) );
fim FAN_N380_7 ( .fault(fault), .net(N380), .FEN(FEN[159]), .op(N380_t7) );
fim FAN_N380_8 ( .fault(fault), .net(N380), .FEN(FEN[160]), .op(N380_t8) );
fim FAN_N380_9 ( .fault(fault), .net(N380), .FEN(FEN[161]), .op(N380_t9) );
fim FAN_N380_10 ( .fault(fault), .net(N380), .FEN(FEN[162]), .op(N380_t10) );
fim FAN_N380_11 ( .fault(fault), .net(N380), .FEN(FEN[163]), .op(N380_t11) );
fim FAN_N393_0 ( .fault(fault), .net(N393), .FEN(FEN[164]), .op(N393_t0) );
fim FAN_N393_1 ( .fault(fault), .net(N393), .FEN(FEN[165]), .op(N393_t1) );
fim FAN_N393_2 ( .fault(fault), .net(N393), .FEN(FEN[166]), .op(N393_t2) );
fim FAN_N393_3 ( .fault(fault), .net(N393), .FEN(FEN[167]), .op(N393_t3) );
fim FAN_N393_4 ( .fault(fault), .net(N393), .FEN(FEN[168]), .op(N393_t4) );
fim FAN_N393_5 ( .fault(fault), .net(N393), .FEN(FEN[169]), .op(N393_t5) );
fim FAN_N393_6 ( .fault(fault), .net(N393), .FEN(FEN[170]), .op(N393_t6) );
fim FAN_N393_7 ( .fault(fault), .net(N393), .FEN(FEN[171]), .op(N393_t7) );
fim FAN_N393_8 ( .fault(fault), .net(N393), .FEN(FEN[172]), .op(N393_t8) );
fim FAN_N393_9 ( .fault(fault), .net(N393), .FEN(FEN[173]), .op(N393_t9) );
fim FAN_N393_10 ( .fault(fault), .net(N393), .FEN(FEN[174]), .op(N393_t10) );
fim FAN_N393_11 ( .fault(fault), .net(N393), .FEN(FEN[175]), .op(N393_t11) );
fim FAN_N419_0 ( .fault(fault), .net(N419), .FEN(FEN[176]), .op(N419_t0) );
fim FAN_N419_1 ( .fault(fault), .net(N419), .FEN(FEN[177]), .op(N419_t1) );
fim FAN_N419_2 ( .fault(fault), .net(N419), .FEN(FEN[178]), .op(N419_t2) );
fim FAN_N419_3 ( .fault(fault), .net(N419), .FEN(FEN[179]), .op(N419_t3) );
fim FAN_N419_4 ( .fault(fault), .net(N419), .FEN(FEN[180]), .op(N419_t4) );
fim FAN_N419_5 ( .fault(fault), .net(N419), .FEN(FEN[181]), .op(N419_t5) );
fim FAN_N419_6 ( .fault(fault), .net(N419), .FEN(FEN[182]), .op(N419_t6) );
fim FAN_N419_7 ( .fault(fault), .net(N419), .FEN(FEN[183]), .op(N419_t7) );
fim FAN_N419_8 ( .fault(fault), .net(N419), .FEN(FEN[184]), .op(N419_t8) );
fim FAN_N419_9 ( .fault(fault), .net(N419), .FEN(FEN[185]), .op(N419_t9) );
fim FAN_N419_10 ( .fault(fault), .net(N419), .FEN(FEN[186]), .op(N419_t10) );
fim FAN_N419_11 ( .fault(fault), .net(N419), .FEN(FEN[187]), .op(N419_t11) );
fim FAN_N445_0 ( .fault(fault), .net(N445), .FEN(FEN[188]), .op(N445_t0) );
fim FAN_N445_1 ( .fault(fault), .net(N445), .FEN(FEN[189]), .op(N445_t1) );
fim FAN_N445_2 ( .fault(fault), .net(N445), .FEN(FEN[190]), .op(N445_t2) );
fim FAN_N445_3 ( .fault(fault), .net(N445), .FEN(FEN[191]), .op(N445_t3) );
fim FAN_N445_4 ( .fault(fault), .net(N445), .FEN(FEN[192]), .op(N445_t4) );
fim FAN_N445_5 ( .fault(fault), .net(N445), .FEN(FEN[193]), .op(N445_t5) );
fim FAN_N445_6 ( .fault(fault), .net(N445), .FEN(FEN[194]), .op(N445_t6) );
fim FAN_N445_7 ( .fault(fault), .net(N445), .FEN(FEN[195]), .op(N445_t7) );
fim FAN_N445_8 ( .fault(fault), .net(N445), .FEN(FEN[196]), .op(N445_t8) );
fim FAN_N445_9 ( .fault(fault), .net(N445), .FEN(FEN[197]), .op(N445_t9) );
fim FAN_N445_10 ( .fault(fault), .net(N445), .FEN(FEN[198]), .op(N445_t10) );
fim FAN_N445_11 ( .fault(fault), .net(N445), .FEN(FEN[199]), .op(N445_t11) );
fim FAN_N432_0 ( .fault(fault), .net(N432), .FEN(FEN[200]), .op(N432_t0) );
fim FAN_N432_1 ( .fault(fault), .net(N432), .FEN(FEN[201]), .op(N432_t1) );
fim FAN_N432_2 ( .fault(fault), .net(N432), .FEN(FEN[202]), .op(N432_t2) );
fim FAN_N432_3 ( .fault(fault), .net(N432), .FEN(FEN[203]), .op(N432_t3) );
fim FAN_N432_4 ( .fault(fault), .net(N432), .FEN(FEN[204]), .op(N432_t4) );
fim FAN_N432_5 ( .fault(fault), .net(N432), .FEN(FEN[205]), .op(N432_t5) );
fim FAN_N432_6 ( .fault(fault), .net(N432), .FEN(FEN[206]), .op(N432_t6) );
fim FAN_N432_7 ( .fault(fault), .net(N432), .FEN(FEN[207]), .op(N432_t7) );
fim FAN_N432_8 ( .fault(fault), .net(N432), .FEN(FEN[208]), .op(N432_t8) );
fim FAN_N432_9 ( .fault(fault), .net(N432), .FEN(FEN[209]), .op(N432_t9) );
fim FAN_N432_10 ( .fault(fault), .net(N432), .FEN(FEN[210]), .op(N432_t10) );
fim FAN_N432_11 ( .fault(fault), .net(N432), .FEN(FEN[211]), .op(N432_t11) );
fim FAN_N406_0 ( .fault(fault), .net(N406), .FEN(FEN[212]), .op(N406_t0) );
fim FAN_N406_1 ( .fault(fault), .net(N406), .FEN(FEN[213]), .op(N406_t1) );
fim FAN_N406_2 ( .fault(fault), .net(N406), .FEN(FEN[214]), .op(N406_t2) );
fim FAN_N406_3 ( .fault(fault), .net(N406), .FEN(FEN[215]), .op(N406_t3) );
fim FAN_N406_4 ( .fault(fault), .net(N406), .FEN(FEN[216]), .op(N406_t4) );
fim FAN_N406_5 ( .fault(fault), .net(N406), .FEN(FEN[217]), .op(N406_t5) );
fim FAN_N406_6 ( .fault(fault), .net(N406), .FEN(FEN[218]), .op(N406_t6) );
fim FAN_N406_7 ( .fault(fault), .net(N406), .FEN(FEN[219]), .op(N406_t7) );
fim FAN_N406_8 ( .fault(fault), .net(N406), .FEN(FEN[220]), .op(N406_t8) );
fim FAN_N406_9 ( .fault(fault), .net(N406), .FEN(FEN[221]), .op(N406_t9) );
fim FAN_N406_10 ( .fault(fault), .net(N406), .FEN(FEN[222]), .op(N406_t10) );
fim FAN_N406_11 ( .fault(fault), .net(N406), .FEN(FEN[223]), .op(N406_t11) );
fim FAN_N602_0 ( .fault(fault), .net(N602), .FEN(FEN[224]), .op(N602_t0) );
fim FAN_N602_1 ( .fault(fault), .net(N602), .FEN(FEN[225]), .op(N602_t1) );
fim FAN_N602_2 ( .fault(fault), .net(N602), .FEN(FEN[226]), .op(N602_t2) );
fim FAN_N602_3 ( .fault(fault), .net(N602), .FEN(FEN[227]), .op(N602_t3) );
fim FAN_N607_0 ( .fault(fault), .net(N607), .FEN(FEN[228]), .op(N607_t0) );
fim FAN_N607_1 ( .fault(fault), .net(N607), .FEN(FEN[229]), .op(N607_t1) );
fim FAN_N607_2 ( .fault(fault), .net(N607), .FEN(FEN[230]), .op(N607_t2) );
fim FAN_N607_3 ( .fault(fault), .net(N607), .FEN(FEN[231]), .op(N607_t3) );
fim FAN_N620_0 ( .fault(fault), .net(N620), .FEN(FEN[232]), .op(N620_t0) );
fim FAN_N620_1 ( .fault(fault), .net(N620), .FEN(FEN[233]), .op(N620_t1) );
fim FAN_N620_2 ( .fault(fault), .net(N620), .FEN(FEN[234]), .op(N620_t2) );
fim FAN_N620_3 ( .fault(fault), .net(N620), .FEN(FEN[235]), .op(N620_t3) );
fim FAN_N625_0 ( .fault(fault), .net(N625), .FEN(FEN[236]), .op(N625_t0) );
fim FAN_N625_1 ( .fault(fault), .net(N625), .FEN(FEN[237]), .op(N625_t1) );
fim FAN_N625_2 ( .fault(fault), .net(N625), .FEN(FEN[238]), .op(N625_t2) );
fim FAN_N625_3 ( .fault(fault), .net(N625), .FEN(FEN[239]), .op(N625_t3) );
fim FAN_N630_0 ( .fault(fault), .net(N630), .FEN(FEN[240]), .op(N630_t0) );
fim FAN_N630_1 ( .fault(fault), .net(N630), .FEN(FEN[241]), .op(N630_t1) );
fim FAN_N630_2 ( .fault(fault), .net(N630), .FEN(FEN[242]), .op(N630_t2) );
fim FAN_N630_3 ( .fault(fault), .net(N630), .FEN(FEN[243]), .op(N630_t3) );
fim FAN_N635_0 ( .fault(fault), .net(N635), .FEN(FEN[244]), .op(N635_t0) );
fim FAN_N635_1 ( .fault(fault), .net(N635), .FEN(FEN[245]), .op(N635_t1) );
fim FAN_N635_2 ( .fault(fault), .net(N635), .FEN(FEN[246]), .op(N635_t2) );
fim FAN_N635_3 ( .fault(fault), .net(N635), .FEN(FEN[247]), .op(N635_t3) );
fim FAN_N640_0 ( .fault(fault), .net(N640), .FEN(FEN[248]), .op(N640_t0) );
fim FAN_N640_1 ( .fault(fault), .net(N640), .FEN(FEN[249]), .op(N640_t1) );
fim FAN_N640_2 ( .fault(fault), .net(N640), .FEN(FEN[250]), .op(N640_t2) );
fim FAN_N640_3 ( .fault(fault), .net(N640), .FEN(FEN[251]), .op(N640_t3) );
fim FAN_N645_0 ( .fault(fault), .net(N645), .FEN(FEN[252]), .op(N645_t0) );
fim FAN_N645_1 ( .fault(fault), .net(N645), .FEN(FEN[253]), .op(N645_t1) );
fim FAN_N645_2 ( .fault(fault), .net(N645), .FEN(FEN[254]), .op(N645_t2) );
fim FAN_N645_3 ( .fault(fault), .net(N645), .FEN(FEN[255]), .op(N645_t3) );
fim FAN_N650_0 ( .fault(fault), .net(N650), .FEN(FEN[256]), .op(N650_t0) );
fim FAN_N650_1 ( .fault(fault), .net(N650), .FEN(FEN[257]), .op(N650_t1) );
fim FAN_N650_2 ( .fault(fault), .net(N650), .FEN(FEN[258]), .op(N650_t2) );
fim FAN_N650_3 ( .fault(fault), .net(N650), .FEN(FEN[259]), .op(N650_t3) );
fim FAN_N655_0 ( .fault(fault), .net(N655), .FEN(FEN[260]), .op(N655_t0) );
fim FAN_N655_1 ( .fault(fault), .net(N655), .FEN(FEN[261]), .op(N655_t1) );
fim FAN_N655_2 ( .fault(fault), .net(N655), .FEN(FEN[262]), .op(N655_t2) );
fim FAN_N655_3 ( .fault(fault), .net(N655), .FEN(FEN[263]), .op(N655_t3) );
initial begin
    FEN <= {263'b0, 1'b1};
    fault <= 1'b0;
    END <= 1'b0;
    //$display("FEN = %.0f, F = %b", FEN, fault);
    end
    always @(posedge(clk) or posedge(rst)) begin
    if(rst == 1) begin
        FEN <= {263'b0, 1'b1};
        fault <= 1'b0;
        END <= 1'b0;
    end
    else if(clk == 1 && INC == 1) begin
        if (FEN == {1'b1,263'b0} && fault == 1'b0) begin
            fault <= 1;
        end
        if (FEN == {1'b1,263'b0} && fault == 1'b1) begin
            END <= 1;
            fault <= 1;
        end
        FEN = {FEN[262:0], FEN[263]};
        if (( FEN[133] || FEN[143] || FEN[145] || FEN[157] || FEN[169] || FEN[181] || FEN[193] || FEN[205] || FEN[217]) && fault == 1) FEN = {FEN[262:0], FEN[263]};
    end
    end
    //always @(FEN or fault) $monitor("FEN = %.0f, F = %b", FEN, fault);
// EndFaultModel

//Anchor
xor XOR2_1 (N250, N1_t0, N5_t0);
xor XOR2_2 (N251, N9_t0, N13_t0);
xor XOR2_3 (N252, N17_t0, N21_t0);
xor XOR2_4 (N253, N25_t0, N29_t0);
xor XOR2_5 (N254, N33_t0, N37_t0);
xor XOR2_6 (N255, N41_t0, N45_t0);
xor XOR2_7 (N256, N49_t0, N53_t0);
xor XOR2_8 (N257, N57_t0, N61_t0);
xor XOR2_9 (N258, N65_t0, N69_t0);
xor XOR2_10 (N259, N73_t0, N77_t0);
xor XOR2_11 (N260, N81_t0, N85_t0);
xor XOR2_12 (N261, N89_t0, N93_t0);
xor XOR2_13 (N262, N97_t0, N101_t0);
xor XOR2_14 (N263, N105_t0, N109_t0);
xor XOR2_15 (N264, N113_t0, N117_t0);
xor XOR2_16 (N265, N121_t0, N125_t0);
and AND2_17 (N266, N129_t, N137_t0);
and AND2_18 (N267, N130_t, N137_t1);
and AND2_19 (N268, N131_t, N137_t2);
and AND2_20 (N269, N132_t, N137_t3);
and AND2_21 (N270, N133_t, N137_t4);
and AND2_22 (N271, N134_t, N137_t5);
and AND2_23 (N272, N135_t, N137_t6);
and AND2_24 (N273, N136_t, N137_t7);
xor XOR2_25 (N274, N1_t1, N17_t1);
xor XOR2_26 (N275, N33_t1, N49_t1);
xor XOR2_27 (N276, N5_t1, N21_t1);
xor XOR2_28 (N277, N37_t1, N53_t1);
xor XOR2_29 (N278, N9_t1, N25_t1);
xor XOR2_30 (N279, N41_t1, N57_t1);
xor XOR2_31 (N280, N13_t1, N29_t1);
xor XOR2_32 (N281, N45_t1, N61_t1);
xor XOR2_33 (N282, N65_t1, N81_t1);
xor XOR2_34 (N283, N97_t1, N113_t1);
xor XOR2_35 (N284, N69_t1, N85_t1);
xor XOR2_36 (N285, N101_t1, N117_t1);
xor XOR2_37 (N286, N73_t1, N89_t1);
xor XOR2_38 (N287, N105_t1, N121_t1);
xor XOR2_39 (N288, N77_t1, N93_t1);
xor XOR2_40 (N289, N109_t1, N125_t1);
xor XOR2_41 (N290, N250, N251);
xor XOR2_42 (N293, N252, N253);
xor XOR2_43 (N296, N254, N255);
xor XOR2_44 (N299, N256, N257);
xor XOR2_45 (N302, N258, N259);
xor XOR2_46 (N305, N260, N261);
xor XOR2_47 (N308, N262, N263);
xor XOR2_48 (N311, N264, N265);
xor XOR2_49 (N314, N274, N275);
xor XOR2_50 (N315, N276, N277);
xor XOR2_51 (N316, N278, N279);
xor XOR2_52 (N317, N280, N281);
xor XOR2_53 (N318, N282, N283);
xor XOR2_54 (N319, N284, N285);
xor XOR2_55 (N320, N286, N287);
xor XOR2_56 (N321, N288, N289);
xor XOR2_57 (N338, N290_t0, N293_t0);
xor XOR2_58 (N339, N296_t0, N299_t0);
xor XOR2_59 (N340, N290_t1, N296_t1);
xor XOR2_60 (N341, N293_t1, N299_t1);
xor XOR2_61 (N342, N302_t0, N305_t0);
xor XOR2_62 (N343, N308_t0, N311_t0);
xor XOR2_63 (N344, N302_t1, N308_t1);
xor XOR2_64 (N345, N305_t1, N311_t1);
xor XOR2_65 (N346, N266, N342);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
xor XOR2_68 (N349, N269, N345);
xor XOR2_69 (N350, N270, N338);
xor XOR2_70 (N351, N271, N339);
xor XOR2_71 (N352, N272, N340);
xor XOR2_72 (N353, N273, N341);
xor XOR2_73 (N354, N314, N346);
xor XOR2_74 (N367, N315, N347);
xor XOR2_75 (N380, N316, N348);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
xor XOR2_78 (N419, N319, N351);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354_t0);
not NOT1_82 (N555, N367_t0);
not NOT1_83 (N556, N380_t0);
not NOT1_84 (N557, N354_t1);
not NOT1_85 (N558, N367_t1);
not NOT1_86 (N559, N393_t0);
not NOT1_87 (N560, N354_t2);
not NOT1_88 (N561, N380_t1);
not NOT1_89 (N562, N393_t1);
not NOT1_90 (N563, N367_t2);
not NOT1_91 (N564, N380_t2);
not NOT1_92 (N565, N393_t2);
not NOT1_93 (N566, N419_t0);
not NOT1_94 (N567, N445_t0);
not NOT1_95 (N568, N419_t1);
not NOT1_96 (N569, N432_t0);
not NOT1_97 (N570, N406_t0);
not NOT1_98 (N571, N445_t1);
not NOT1_99 (N572, N406_t1);
not NOT1_100 (N573, N432_t1);
not NOT1_101 (N574, N406_t2);
not NOT1_102 (N575, N419_t2);
not NOT1_103 (N576, N432_t2);
not NOT1_104 (N577, N406_t3);
not NOT1_105 (N578, N419_t3);
not NOT1_106 (N579, N445_t2);
not NOT1_107 (N580, N406_t4);
not NOT1_108 (N581, N432_t3);
not NOT1_109 (N582, N445_t3);
not NOT1_110 (N583, N419_t4);
not NOT1_111 (N584, N432_t4);
not NOT1_112 (N585, N445_t4);
not NOT1_113 (N586, N367_t3);
not NOT1_114 (N587, N393_t3);
not NOT1_115 (N588, N367_t4);
not NOT1_116 (N589, N380_t3);
not NOT1_117 (N590, N354_t3);
not NOT1_118 (N591, N393_t4);
not NOT1_119 (N592, N354_t4);
not NOT1_120 (N593, N380_t4);
and AND4_121 (N594, N554, N555, N556, N393_t5);
and AND4_122 (N595, N557, N558, N380_t5, N559);
and AND4_123 (N596, N560, N367_t5, N561, N562);
and AND4_124 (N597, N354_t5, N563, N564, N565);
and AND4_125 (N598, N574, N575, N576, N445_t5);
and AND4_126 (N599, N577, N578, N432_t5, N579);
and AND4_127 (N600, N580, N419_t5, N581, N582);
and AND4_128 (N601, N406_t5, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
or OR4_130 (N607, N598, N599, N600, N601);
and AND5_131 (N620, N406_t6, N566, N432_t6, N567, N602_t0);
and AND5_132 (N625, N406_t7, N568, N569, N445_t6, N602_t1);
and AND5_133 (N630, N570, N419_t6, N432_t7, N571, N602_t2);
and AND5_134 (N635, N572, N419_t7, N573, N445_t7, N602_t3);
and AND5_135 (N640, N354_t6, N586, N380_t6, N587, N607_t0);
and AND5_136 (N645, N354_t7, N588, N589, N393_t6, N607_t1);
and AND5_137 (N650, N590, N367_t6, N380_t7, N591, N607_t2);
and AND5_138 (N655, N592, N367_t7, N593, N393_t7, N607_t3);
and AND2_139 (N692, N354_t8, N620_t0);
and AND2_140 (N693, N367_t8, N620_t1);
and AND2_141 (N694, N380_t8, N620_t2);
and AND2_142 (N695, N393_t8, N620_t3);
and AND2_143 (N696, N354_t9, N625_t0);
and AND2_144 (N697, N367_t9, N625_t1);
and AND2_145 (N698, N380_t9, N625_t2);
and AND2_146 (N699, N393_t9, N625_t3);
and AND2_147 (N700, N354_t10, N630_t0);
and AND2_148 (N701, N367_t10, N630_t1);
and AND2_149 (N702, N380_t10, N630_t2);
and AND2_150 (N703, N393_t10, N630_t3);
and AND2_151 (N704, N354_t11, N635_t0);
and AND2_152 (N705, N367_t11, N635_t1);
and AND2_153 (N706, N380_t11, N635_t2);
and AND2_154 (N707, N393_t11, N635_t3);
and AND2_155 (N708, N406_t8, N640_t0);
and AND2_156 (N709, N419_t8, N640_t1);
and AND2_157 (N710, N432_t8, N640_t2);
and AND2_158 (N711, N445_t8, N640_t3);
and AND2_159 (N712, N406_t9, N645_t0);
and AND2_160 (N713, N419_t9, N645_t1);
and AND2_161 (N714, N432_t9, N645_t2);
and AND2_162 (N715, N445_t9, N645_t3);
and AND2_163 (N716, N406_t10, N650_t0);
and AND2_164 (N717, N419_t10, N650_t1);
and AND2_165 (N718, N432_t10, N650_t2);
and AND2_166 (N719, N445_t10, N650_t3);
and AND2_167 (N720, N406_t11, N655_t0);
and AND2_168 (N721, N419_t11, N655_t1);
and AND2_169 (N722, N432_t11, N655_t2);
and AND2_170 (N723, N445_t11, N655_t3);
xor XOR2_171 (N724, N1_t2, N692);
xor XOR2_172 (N725, N5_t2, N693);
xor XOR2_173 (N726, N9_t2, N694);
xor XOR2_174 (N727, N13_t2, N695);
xor XOR2_175 (N728, N17_t2, N696);
xor XOR2_176 (N729, N21_t2, N697);
xor XOR2_177 (N730, N25_t2, N698);
xor XOR2_178 (N731, N29_t2, N699);
xor XOR2_179 (N732, N33_t2, N700);
xor XOR2_180 (N733, N37_t2, N701);
xor XOR2_181 (N734, N41_t2, N702);
xor XOR2_182 (N735, N45_t2, N703);
xor XOR2_183 (N736, N49_t2, N704);
xor XOR2_184 (N737, N53_t2, N705);
xor XOR2_185 (N738, N57_t2, N706);
xor XOR2_186 (N739, N61_t2, N707);
xor XOR2_187 (N740, N65_t2, N708);
xor XOR2_188 (N741, N69_t2, N709);
xor XOR2_189 (N742, N73_t2, N710);
xor XOR2_190 (N743, N77_t2, N711);
xor XOR2_191 (N744, N81_t2, N712);
xor XOR2_192 (N745, N85_t2, N713);
xor XOR2_193 (N746, N89_t2, N714);
xor XOR2_194 (N747, N93_t2, N715);
xor XOR2_195 (N748, N97_t2, N716);
xor XOR2_196 (N749, N101_t2, N717);
xor XOR2_197 (N750, N105_t2, N718);
xor XOR2_198 (N751, N109_t2, N719);
xor XOR2_199 (N752, N113_t2, N720);
xor XOR2_200 (N753, N117_t2, N721);
xor XOR2_201 (N754, N121_t2, N722);
xor XOR2_202 (N755, N125_t2, N723);

endmodule
